//Generate the verilog at 2025-02-27T22:05:00
module Top (
clock,
io_clrn,
io_ps2_clk,
io_ps2_data,
reset,
io_seg_out_0,
io_seg_out_1,
io_seg_out_2,
io_seg_out_3,
io_seg_out_4,
io_seg_out_5
);

input clock ;
input io_clrn ;
input io_ps2_clk ;
input io_ps2_data ;
input reset ;
output [7:0] io_seg_out_0 ;
output [7:0] io_seg_out_1 ;
output [7:0] io_seg_out_2 ;
output [7:0] io_seg_out_3 ;
output [7:0] io_seg_out_4 ;
output [7:0] io_seg_out_5 ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire counter_io_key_press ;
wire counter_io_key_release ;
wire display_en ;
wire keyboard_io_nextdata_n ;
wire keyboard_io_ready ;
wire ready_delay ;
wire \counter/_000_ ;
wire \counter/_001_ ;
wire \counter/_002_ ;
wire \counter/_003_ ;
wire \counter/_004_ ;
wire \counter/_005_ ;
wire \counter/_006_ ;
wire \counter/_007_ ;
wire \counter/_008_ ;
wire \counter/_009_ ;
wire \counter/_010_ ;
wire \counter/_011_ ;
wire \counter/_012_ ;
wire \counter/_013_ ;
wire \counter/_014_ ;
wire \counter/_015_ ;
wire \counter/_016_ ;
wire \counter/_017_ ;
wire \counter/_018_ ;
wire \counter/_019_ ;
wire \counter/_020_ ;
wire \counter/_021_ ;
wire \counter/_022_ ;
wire \counter/_023_ ;
wire \counter/_024_ ;
wire \counter/_025_ ;
wire \counter/_026_ ;
wire \counter/_027_ ;
wire \counter/_028_ ;
wire \counter/_029_ ;
wire \counter/_030_ ;
wire \counter/_031_ ;
wire \counter/_032_ ;
wire \counter/_033_ ;
wire \counter/_034_ ;
wire \counter/_035_ ;
wire \counter/_036_ ;
wire \counter/_037_ ;
wire \counter/_038_ ;
wire \counter/_039_ ;
wire \counter/_040_ ;
wire \counter/_041_ ;
wire \counter/_042_ ;
wire \counter/_043_ ;
wire \counter/_044_ ;
wire \counter/_045_ ;
wire \counter/_046_ ;
wire \counter/_047_ ;
wire \counter/_048_ ;
wire \counter/_049_ ;
wire \counter/_050_ ;
wire \counter/_051_ ;
wire \counter/_052_ ;
wire \counter/_053_ ;
wire \counter/_054_ ;
wire \counter/_055_ ;
wire \counter/_056_ ;
wire \counter/_057_ ;
wire \counter/_058_ ;
wire \counter/_059_ ;
wire \counter/_060_ ;
wire \counter/_061_ ;
wire \counter/_062_ ;
wire \counter/_063_ ;
wire \counter/_064_ ;
wire \counter/_065_ ;
wire \counter/_066_ ;
wire \counter/_067_ ;
wire \counter/_068_ ;
wire \counter/_069_ ;
wire \counter/_070_ ;
wire \counter/_071_ ;
wire \counter/_072_ ;
wire \counter/_073_ ;
wire \counter/_074_ ;
wire \counter/_075_ ;
wire \counter/_076_ ;
wire \counter/_077_ ;
wire \counter/_078_ ;
wire \counter/_079_ ;
wire \counter/_080_ ;
wire \counter/_081_ ;
wire \counter/_082_ ;
wire \counter/_083_ ;
wire \counter/counted ;
wire \decoder/_000_ ;
wire \decoder/_001_ ;
wire \decoder/_002_ ;
wire \decoder/_003_ ;
wire \decoder/_004_ ;
wire \decoder/_005_ ;
wire \decoder/_006_ ;
wire \decoder/_007_ ;
wire \decoder/_008_ ;
wire \decoder/_009_ ;
wire \decoder/_010_ ;
wire \decoder/_011_ ;
wire \decoder/_012_ ;
wire \decoder/_013_ ;
wire \decoder/_014_ ;
wire \decoder/_015_ ;
wire \decoder/_016_ ;
wire \decoder/_017_ ;
wire \decoder/_018_ ;
wire \decoder/_019_ ;
wire \decoder/_020_ ;
wire \decoder/_021_ ;
wire \decoder/_022_ ;
wire \decoder/_023_ ;
wire \decoder/_024_ ;
wire \decoder/_025_ ;
wire \decoder/_026_ ;
wire \decoder/_027_ ;
wire \decoder/_028_ ;
wire \decoder/_029_ ;
wire \decoder/_030_ ;
wire \decoder/_031_ ;
wire \decoder/_032_ ;
wire \decoder/_033_ ;
wire \decoder/_034_ ;
wire \decoder/_035_ ;
wire \decoder/_036_ ;
wire \decoder/_037_ ;
wire \decoder/_038_ ;
wire \decoder/_039_ ;
wire \decoder/_040_ ;
wire \decoder/_041_ ;
wire \decoder/_042_ ;
wire \decoder/_043_ ;
wire \decoder/_044_ ;
wire \decoder/_045_ ;
wire \decoder/_046_ ;
wire \decoder/_047_ ;
wire \decoder/_048_ ;
wire \decoder/_049_ ;
wire \decoder/_050_ ;
wire \decoder/_051_ ;
wire \decoder/_052_ ;
wire \decoder/_053_ ;
wire \decoder/_054_ ;
wire \decoder/_055_ ;
wire \decoder/_056_ ;
wire \decoder/_057_ ;
wire \decoder/_058_ ;
wire \decoder/_059_ ;
wire \decoder/_060_ ;
wire \decoder/_061_ ;
wire \decoder/_062_ ;
wire \decoder/_063_ ;
wire \decoder/_064_ ;
wire \decoder/_065_ ;
wire \decoder/_066_ ;
wire \decoder/_067_ ;
wire \decoder/_068_ ;
wire \decoder/_069_ ;
wire \decoder/_070_ ;
wire \decoder/_071_ ;
wire \decoder/_072_ ;
wire \decoder/_073_ ;
wire \decoder/_074_ ;
wire \decoder/_075_ ;
wire \decoder/_076_ ;
wire \decoder/_077_ ;
wire \decoder/_078_ ;
wire \decoder/_079_ ;
wire \decoder/_080_ ;
wire \decoder/_081_ ;
wire \decoder/_082_ ;
wire \decoder/_083_ ;
wire \decoder/_084_ ;
wire \decoder/_085_ ;
wire \decoder/_086_ ;
wire \decoder/_087_ ;
wire \decoder/_088_ ;
wire \decoder/_089_ ;
wire \decoder/_090_ ;
wire \decoder/_091_ ;
wire \decoder/_092_ ;
wire \decoder/_093_ ;
wire \decoder/_094_ ;
wire \decoder/_095_ ;
wire \decoder/_096_ ;
wire \decoder/_097_ ;
wire \decoder/_098_ ;
wire \decoder/_099_ ;
wire \decoder/_100_ ;
wire \decoder/_101_ ;
wire \decoder/_102_ ;
wire \decoder/_103_ ;
wire \decoder/_104_ ;
wire \decoder/_105_ ;
wire \decoder/_106_ ;
wire \decoder/_107_ ;
wire \decoder/_108_ ;
wire \decoder/_109_ ;
wire \decoder/_110_ ;
wire \decoder/_111_ ;
wire \decoder/_112_ ;
wire \decoder/_113_ ;
wire \decoder/_114_ ;
wire \decoder/_115_ ;
wire \decoder/_116_ ;
wire \decoder/_117_ ;
wire \decoder/_118_ ;
wire \decoder/_119_ ;
wire \decoder/_120_ ;
wire \decoder/_121_ ;
wire \decoder/_122_ ;
wire \decoder/_123_ ;
wire \decoder/_124_ ;
wire \decoder/_125_ ;
wire \decoder/_126_ ;
wire \decoder/_127_ ;
wire \decoder/_128_ ;
wire \decoder/_129_ ;
wire \decoder/_130_ ;
wire \decoder/_131_ ;
wire \decoder/_132_ ;
wire \decoder/isBreakCode ;
wire \keyboard/_0000_ ;
wire \keyboard/_0001_ ;
wire \keyboard/_0002_ ;
wire \keyboard/_0003_ ;
wire \keyboard/_0004_ ;
wire \keyboard/_0005_ ;
wire \keyboard/_0006_ ;
wire \keyboard/_0007_ ;
wire \keyboard/_0008_ ;
wire \keyboard/_0009_ ;
wire \keyboard/_0010_ ;
wire \keyboard/_0011_ ;
wire \keyboard/_0012_ ;
wire \keyboard/_0013_ ;
wire \keyboard/_0014_ ;
wire \keyboard/_0015_ ;
wire \keyboard/_0016_ ;
wire \keyboard/_0017_ ;
wire \keyboard/_0018_ ;
wire \keyboard/_0019_ ;
wire \keyboard/_0020_ ;
wire \keyboard/_0021_ ;
wire \keyboard/_0022_ ;
wire \keyboard/_0023_ ;
wire \keyboard/_0024_ ;
wire \keyboard/_0025_ ;
wire \keyboard/_0026_ ;
wire \keyboard/_0027_ ;
wire \keyboard/_0028_ ;
wire \keyboard/_0029_ ;
wire \keyboard/_0030_ ;
wire \keyboard/_0031_ ;
wire \keyboard/_0032_ ;
wire \keyboard/_0033_ ;
wire \keyboard/_0034_ ;
wire \keyboard/_0035_ ;
wire \keyboard/_0036_ ;
wire \keyboard/_0037_ ;
wire \keyboard/_0038_ ;
wire \keyboard/_0039_ ;
wire \keyboard/_0040_ ;
wire \keyboard/_0041_ ;
wire \keyboard/_0042_ ;
wire \keyboard/_0043_ ;
wire \keyboard/_0044_ ;
wire \keyboard/_0045_ ;
wire \keyboard/_0046_ ;
wire \keyboard/_0047_ ;
wire \keyboard/_0048_ ;
wire \keyboard/_0049_ ;
wire \keyboard/_0050_ ;
wire \keyboard/_0051_ ;
wire \keyboard/_0052_ ;
wire \keyboard/_0053_ ;
wire \keyboard/_0054_ ;
wire \keyboard/_0055_ ;
wire \keyboard/_0056_ ;
wire \keyboard/_0057_ ;
wire \keyboard/_0058_ ;
wire \keyboard/_0059_ ;
wire \keyboard/_0060_ ;
wire \keyboard/_0061_ ;
wire \keyboard/_0062_ ;
wire \keyboard/_0063_ ;
wire \keyboard/_0064_ ;
wire \keyboard/_0065_ ;
wire \keyboard/_0066_ ;
wire \keyboard/_0067_ ;
wire \keyboard/_0068_ ;
wire \keyboard/_0069_ ;
wire \keyboard/_0070_ ;
wire \keyboard/_0071_ ;
wire \keyboard/_0072_ ;
wire \keyboard/_0073_ ;
wire \keyboard/_0074_ ;
wire \keyboard/_0075_ ;
wire \keyboard/_0076_ ;
wire \keyboard/_0077_ ;
wire \keyboard/_0078_ ;
wire \keyboard/_0079_ ;
wire \keyboard/_0080_ ;
wire \keyboard/_0081_ ;
wire \keyboard/_0082_ ;
wire \keyboard/_0083_ ;
wire \keyboard/_0084_ ;
wire \keyboard/_0085_ ;
wire \keyboard/_0086_ ;
wire \keyboard/_0087_ ;
wire \keyboard/_0088_ ;
wire \keyboard/_0089_ ;
wire \keyboard/_0090_ ;
wire \keyboard/_0091_ ;
wire \keyboard/_0092_ ;
wire \keyboard/_0093_ ;
wire \keyboard/_0094_ ;
wire \keyboard/_0095_ ;
wire \keyboard/_0096_ ;
wire \keyboard/_0097_ ;
wire \keyboard/_0098_ ;
wire \keyboard/_0099_ ;
wire \keyboard/_0100_ ;
wire \keyboard/_0101_ ;
wire \keyboard/_0102_ ;
wire \keyboard/_0103_ ;
wire \keyboard/_0104_ ;
wire \keyboard/_0105_ ;
wire \keyboard/_0106_ ;
wire \keyboard/_0107_ ;
wire \keyboard/_0108_ ;
wire \keyboard/_0109_ ;
wire \keyboard/_0110_ ;
wire \keyboard/_0111_ ;
wire \keyboard/_0112_ ;
wire \keyboard/_0113_ ;
wire \keyboard/_0114_ ;
wire \keyboard/_0115_ ;
wire \keyboard/_0116_ ;
wire \keyboard/_0117_ ;
wire \keyboard/_0118_ ;
wire \keyboard/_0119_ ;
wire \keyboard/_0120_ ;
wire \keyboard/_0121_ ;
wire \keyboard/_0122_ ;
wire \keyboard/_0123_ ;
wire \keyboard/_0124_ ;
wire \keyboard/_0125_ ;
wire \keyboard/_0126_ ;
wire \keyboard/_0127_ ;
wire \keyboard/_0128_ ;
wire \keyboard/_0129_ ;
wire \keyboard/_0130_ ;
wire \keyboard/_0131_ ;
wire \keyboard/_0132_ ;
wire \keyboard/_0133_ ;
wire \keyboard/_0134_ ;
wire \keyboard/_0135_ ;
wire \keyboard/_0136_ ;
wire \keyboard/_0137_ ;
wire \keyboard/_0138_ ;
wire \keyboard/_0139_ ;
wire \keyboard/_0140_ ;
wire \keyboard/_0141_ ;
wire \keyboard/_0142_ ;
wire \keyboard/_0143_ ;
wire \keyboard/_0144_ ;
wire \keyboard/_0145_ ;
wire \keyboard/_0146_ ;
wire \keyboard/_0147_ ;
wire \keyboard/_0148_ ;
wire \keyboard/_0149_ ;
wire \keyboard/_0150_ ;
wire \keyboard/_0151_ ;
wire \keyboard/_0152_ ;
wire \keyboard/_0153_ ;
wire \keyboard/_0154_ ;
wire \keyboard/_0155_ ;
wire \keyboard/_0156_ ;
wire \keyboard/_0157_ ;
wire \keyboard/_0158_ ;
wire \keyboard/_0159_ ;
wire \keyboard/_0160_ ;
wire \keyboard/_0161_ ;
wire \keyboard/_0162_ ;
wire \keyboard/_0163_ ;
wire \keyboard/_0164_ ;
wire \keyboard/_0165_ ;
wire \keyboard/_0166_ ;
wire \keyboard/_0167_ ;
wire \keyboard/_0168_ ;
wire \keyboard/_0169_ ;
wire \keyboard/_0170_ ;
wire \keyboard/_0171_ ;
wire \keyboard/_0172_ ;
wire \keyboard/_0173_ ;
wire \keyboard/_0174_ ;
wire \keyboard/_0175_ ;
wire \keyboard/_0176_ ;
wire \keyboard/_0177_ ;
wire \keyboard/_0178_ ;
wire \keyboard/_0179_ ;
wire \keyboard/_0180_ ;
wire \keyboard/_0181_ ;
wire \keyboard/_0182_ ;
wire \keyboard/_0183_ ;
wire \keyboard/_0184_ ;
wire \keyboard/_0185_ ;
wire \keyboard/_0186_ ;
wire \keyboard/_0187_ ;
wire \keyboard/_0188_ ;
wire \keyboard/_0189_ ;
wire \keyboard/_0190_ ;
wire \keyboard/_0191_ ;
wire \keyboard/_0192_ ;
wire \keyboard/_0193_ ;
wire \keyboard/_0194_ ;
wire \keyboard/_0195_ ;
wire \keyboard/_0196_ ;
wire \keyboard/_0197_ ;
wire \keyboard/_0198_ ;
wire \keyboard/_0199_ ;
wire \keyboard/_0200_ ;
wire \keyboard/_0201_ ;
wire \keyboard/_0202_ ;
wire \keyboard/_0203_ ;
wire \keyboard/_0204_ ;
wire \keyboard/_0205_ ;
wire \keyboard/_0206_ ;
wire \keyboard/_0207_ ;
wire \keyboard/_0208_ ;
wire \keyboard/_0209_ ;
wire \keyboard/_0210_ ;
wire \keyboard/_0211_ ;
wire \keyboard/_0212_ ;
wire \keyboard/_0213_ ;
wire \keyboard/_0214_ ;
wire \keyboard/_0215_ ;
wire \keyboard/_0216_ ;
wire \keyboard/_0217_ ;
wire \keyboard/_0218_ ;
wire \keyboard/_0219_ ;
wire \keyboard/_0220_ ;
wire \keyboard/_0221_ ;
wire \keyboard/_0222_ ;
wire \keyboard/_0223_ ;
wire \keyboard/_0224_ ;
wire \keyboard/_0225_ ;
wire \keyboard/_0226_ ;
wire \keyboard/_0227_ ;
wire \keyboard/_0228_ ;
wire \keyboard/_0229_ ;
wire \keyboard/_0230_ ;
wire \keyboard/_0231_ ;
wire \keyboard/_0232_ ;
wire \keyboard/_0233_ ;
wire \keyboard/_0234_ ;
wire \keyboard/_0235_ ;
wire \keyboard/_0236_ ;
wire \keyboard/_0237_ ;
wire \keyboard/_0238_ ;
wire \keyboard/_0239_ ;
wire \keyboard/_0240_ ;
wire \keyboard/_0241_ ;
wire \keyboard/_0242_ ;
wire \keyboard/_0243_ ;
wire \keyboard/_0244_ ;
wire \keyboard/_0245_ ;
wire \keyboard/_0246_ ;
wire \keyboard/_0247_ ;
wire \keyboard/_0248_ ;
wire \keyboard/_0249_ ;
wire \keyboard/_0250_ ;
wire \keyboard/_0251_ ;
wire \keyboard/_0252_ ;
wire \keyboard/_0253_ ;
wire \keyboard/_0254_ ;
wire \keyboard/_0255_ ;
wire \keyboard/_0256_ ;
wire \keyboard/_0257_ ;
wire \keyboard/_0258_ ;
wire \keyboard/_0259_ ;
wire \keyboard/_0260_ ;
wire \keyboard/_0261_ ;
wire \keyboard/_0262_ ;
wire \keyboard/_0263_ ;
wire \keyboard/_0264_ ;
wire \keyboard/_0265_ ;
wire \keyboard/_0266_ ;
wire \keyboard/_0267_ ;
wire \keyboard/_0268_ ;
wire \keyboard/_0269_ ;
wire \keyboard/_0270_ ;
wire \keyboard/_0271_ ;
wire \keyboard/_0272_ ;
wire \keyboard/_0273_ ;
wire \keyboard/_0274_ ;
wire \keyboard/_0275_ ;
wire \keyboard/_0276_ ;
wire \keyboard/_0277_ ;
wire \keyboard/_0278_ ;
wire \keyboard/_0279_ ;
wire \keyboard/_0280_ ;
wire \keyboard/_0281_ ;
wire \keyboard/_0282_ ;
wire \keyboard/_0283_ ;
wire \keyboard/_0284_ ;
wire \keyboard/_0285_ ;
wire \keyboard/_0286_ ;
wire \keyboard/_0287_ ;
wire \keyboard/_0288_ ;
wire \keyboard/_0289_ ;
wire \keyboard/_0290_ ;
wire \keyboard/_0291_ ;
wire \keyboard/_0292_ ;
wire \keyboard/_0293_ ;
wire \keyboard/_0294_ ;
wire \keyboard/_0295_ ;
wire \keyboard/_0296_ ;
wire \keyboard/_0297_ ;
wire \keyboard/_0298_ ;
wire \keyboard/_0299_ ;
wire \keyboard/_0300_ ;
wire \keyboard/_0301_ ;
wire \keyboard/_0302_ ;
wire \keyboard/_0303_ ;
wire \keyboard/_0304_ ;
wire \keyboard/_0305_ ;
wire \keyboard/_0306_ ;
wire \keyboard/_0307_ ;
wire \keyboard/_0308_ ;
wire \keyboard/_0309_ ;
wire \keyboard/_0310_ ;
wire \keyboard/_0311_ ;
wire \keyboard/_0312_ ;
wire \keyboard/_0313_ ;
wire \keyboard/_0314_ ;
wire \keyboard/_0315_ ;
wire \keyboard/_0316_ ;
wire \keyboard/_0317_ ;
wire \keyboard/_0318_ ;
wire \keyboard/_0319_ ;
wire \keyboard/_0320_ ;
wire \keyboard/_0321_ ;
wire \keyboard/_0322_ ;
wire \keyboard/_0323_ ;
wire \keyboard/_0324_ ;
wire \keyboard/_0325_ ;
wire \keyboard/_0326_ ;
wire \keyboard/_0327_ ;
wire \keyboard/_0328_ ;
wire \keyboard/_0329_ ;
wire \keyboard/_0330_ ;
wire \keyboard/_0331_ ;
wire \keyboard/_0332_ ;
wire \keyboard/_0333_ ;
wire \keyboard/_0334_ ;
wire \keyboard/_0335_ ;
wire \keyboard/_0336_ ;
wire \keyboard/_0337_ ;
wire \keyboard/_0338_ ;
wire \keyboard/_0339_ ;
wire \keyboard/_0340_ ;
wire \keyboard/_0341_ ;
wire \keyboard/_0342_ ;
wire \keyboard/_0343_ ;
wire \keyboard/_0344_ ;
wire \keyboard/_0345_ ;
wire \keyboard/_0346_ ;
wire \keyboard/_0347_ ;
wire \keyboard/_0348_ ;
wire \keyboard/_0349_ ;
wire \keyboard/_0350_ ;
wire \keyboard/_0351_ ;
wire \keyboard/_0352_ ;
wire \keyboard/_0353_ ;
wire \keyboard/_0354_ ;
wire \keyboard/_0355_ ;
wire \keyboard/_0356_ ;
wire \keyboard/_0357_ ;
wire \keyboard/_0358_ ;
wire \keyboard/_0359_ ;
wire \keyboard/_0360_ ;
wire \keyboard/_0361_ ;
wire \keyboard/_0362_ ;
wire \keyboard/_0363_ ;
wire \keyboard/_0364_ ;
wire \keyboard/_0365_ ;
wire \keyboard/_0366_ ;
wire \keyboard/_0367_ ;
wire \keyboard/_0368_ ;
wire \keyboard/_0369_ ;
wire \keyboard/_0370_ ;
wire \keyboard/_0371_ ;
wire \keyboard/_0372_ ;
wire \keyboard/_0373_ ;
wire \keyboard/_0374_ ;
wire \keyboard/_0375_ ;
wire \keyboard/_0376_ ;
wire \keyboard/_0377_ ;
wire \keyboard/_0378_ ;
wire \keyboard/_0379_ ;
wire \keyboard/_0380_ ;
wire \keyboard/_0381_ ;
wire \keyboard/_0382_ ;
wire \keyboard/_0383_ ;
wire \keyboard/_0384_ ;
wire \keyboard/_0385_ ;
wire \keyboard/_0386_ ;
wire \keyboard/_0387_ ;
wire \keyboard/_0388_ ;
wire \keyboard/_0389_ ;
wire \keyboard/_0390_ ;
wire \keyboard/_0391_ ;
wire \keyboard/_0392_ ;
wire \keyboard/_0393_ ;
wire \keyboard/_0394_ ;
wire \keyboard/_0395_ ;
wire \keyboard/_0396_ ;
wire \keyboard/_0397_ ;
wire \keyboard/_0398_ ;
wire \keyboard/_0399_ ;
wire \keyboard/_0400_ ;
wire \keyboard/_0401_ ;
wire \keyboard/_0402_ ;
wire \keyboard/_0403_ ;
wire \keyboard/_0404_ ;
wire \keyboard/_0405_ ;
wire \keyboard/_0406_ ;
wire \keyboard/_0407_ ;
wire \keyboard/_0408_ ;
wire \keyboard/_0409_ ;
wire \keyboard/_0410_ ;
wire \keyboard/_0411_ ;
wire \keyboard/_0412_ ;
wire \keyboard/_0413_ ;
wire \keyboard/_0414_ ;
wire \keyboard/_0415_ ;
wire \keyboard/_0416_ ;
wire \keyboard/_0417_ ;
wire \keyboard/_0418_ ;
wire \keyboard/_0419_ ;
wire \keyboard/_0420_ ;
wire \keyboard/_0421_ ;
wire \keyboard/_0422_ ;
wire \keyboard/_0423_ ;
wire \keyboard/_0424_ ;
wire \keyboard/_0425_ ;
wire \keyboard/_0426_ ;
wire \keyboard/_0427_ ;
wire \keyboard/_0428_ ;
wire \keyboard/_0429_ ;
wire \keyboard/_0430_ ;
wire \keyboard/_0431_ ;
wire \keyboard/_0432_ ;
wire \keyboard/_0433_ ;
wire \keyboard/_0434_ ;
wire \keyboard/_0435_ ;
wire \keyboard/_0436_ ;
wire \keyboard/_0437_ ;
wire \keyboard/_0438_ ;
wire \keyboard/_0439_ ;
wire \keyboard/_0440_ ;
wire \keyboard/_0441_ ;
wire \keyboard/_0442_ ;
wire \keyboard/_0443_ ;
wire \keyboard/_0444_ ;
wire \keyboard/_0445_ ;
wire \keyboard/_0446_ ;
wire \keyboard/_0447_ ;
wire \keyboard/_0448_ ;
wire \keyboard/_0449_ ;
wire \keyboard/_0450_ ;
wire \keyboard/_0451_ ;
wire \keyboard/_0452_ ;
wire \keyboard/_0453_ ;
wire \keyboard/_0454_ ;
wire \keyboard/_0455_ ;
wire \keyboard/_0456_ ;
wire \keyboard/_0457_ ;
wire \keyboard/_0458_ ;
wire \keyboard/_0459_ ;
wire \keyboard/_0460_ ;
wire \keyboard/_0461_ ;
wire \keyboard/_0462_ ;
wire \keyboard/_0463_ ;
wire \keyboard/_0464_ ;
wire \keyboard/_0465_ ;
wire \keyboard/_0466_ ;
wire \keyboard/_0467_ ;
wire \keyboard/_0468_ ;
wire \keyboard/_0469_ ;
wire \keyboard/_0470_ ;
wire \keyboard/_0471_ ;
wire \keyboard/_0472_ ;
wire \keyboard/_0473_ ;
wire \keyboard/_0474_ ;
wire \keyboard/_0475_ ;
wire \keyboard/_0476_ ;
wire \keyboard/_0477_ ;
wire \keyboard/_0478_ ;
wire \keyboard/_0479_ ;
wire \keyboard/_0480_ ;
wire \keyboard/_0481_ ;
wire \keyboard/_0482_ ;
wire \keyboard/_0483_ ;
wire \keyboard/_0484_ ;
wire \keyboard/_0485_ ;
wire \keyboard/_0486_ ;
wire \keyboard/_0487_ ;
wire \keyboard/_0488_ ;
wire \keyboard/_0489_ ;
wire \keyboard/_0490_ ;
wire \keyboard/_0491_ ;
wire \keyboard/_0492_ ;
wire \keyboard/_0493_ ;
wire \keyboard/_0494_ ;
wire \keyboard/_0495_ ;
wire \keyboard/_0496_ ;
wire \keyboard/_0497_ ;
wire \keyboard/_0498_ ;
wire \keyboard/_0499_ ;
wire \keyboard/_0500_ ;
wire \keyboard/_0501_ ;
wire \keyboard/_0502_ ;
wire \keyboard/_0503_ ;
wire \keyboard/_0504_ ;
wire \keyboard/_0505_ ;
wire \keyboard/_0506_ ;
wire \keyboard/_0507_ ;
wire \keyboard/_0508_ ;
wire \keyboard/_0509_ ;
wire \keyboard/_0510_ ;
wire \keyboard/_0511_ ;
wire \keyboard/_0512_ ;
wire \keyboard/_0513_ ;
wire \keyboard/_0514_ ;
wire \keyboard/_0515_ ;
wire \keyboard/_0516_ ;
wire \keyboard/_0517_ ;
wire \keyboard/_0518_ ;
wire \keyboard/_0519_ ;
wire \keyboard/_0520_ ;
wire \keyboard/_0521_ ;
wire \keyboard/_0522_ ;
wire \keyboard/_0523_ ;
wire \keyboard/_0524_ ;
wire \keyboard/_0525_ ;
wire \keyboard/_0526_ ;
wire \keyboard/_0527_ ;
wire \keyboard/_0528_ ;
wire \keyboard/_0529_ ;
wire \keyboard/_0530_ ;
wire \keyboard/_0531_ ;
wire \keyboard/_0532_ ;
wire \keyboard/_0533_ ;
wire \keyboard/_0534_ ;
wire \keyboard/_0535_ ;
wire \keyboard/_0536_ ;
wire \keyboard/_0537_ ;
wire \keyboard/_0538_ ;
wire \keyboard/_0539_ ;
wire \keyboard/_0540_ ;
wire \keyboard/_0541_ ;
wire \keyboard/_0542_ ;
wire \keyboard/_0543_ ;
wire \keyboard/_0544_ ;
wire \keyboard/_0545_ ;
wire \keyboard/_0546_ ;
wire \keyboard/_0547_ ;
wire \keyboard/_0548_ ;
wire \keyboard/_0549_ ;
wire \keyboard/_0550_ ;
wire \keyboard/_0551_ ;
wire \keyboard/_0552_ ;
wire \keyboard/_0553_ ;
wire \keyboard/_0554_ ;
wire \keyboard/_0555_ ;
wire \keyboard/_0556_ ;
wire \keyboard/_0557_ ;
wire \keyboard/_0558_ ;
wire \keyboard/_0559_ ;
wire \keyboard/_0560_ ;
wire \keyboard/_0561_ ;
wire \keyboard/_0562_ ;
wire \keyboard/_0563_ ;
wire \keyboard/_0564_ ;
wire \keyboard/_0565_ ;
wire \keyboard/_0566_ ;
wire \keyboard/_0567_ ;
wire \keyboard/_0568_ ;
wire \keyboard/_0569_ ;
wire \keyboard/_0570_ ;
wire \keyboard/_0571_ ;
wire \keyboard/_0572_ ;
wire \keyboard/_0573_ ;
wire \keyboard/_0574_ ;
wire \keyboard/_0575_ ;
wire \keyboard/_0576_ ;
wire \keyboard/_0577_ ;
wire \keyboard/_0578_ ;
wire \keyboard/_0579_ ;
wire \keyboard/_0580_ ;
wire \keyboard/_0581_ ;
wire \keyboard/_0582_ ;
wire \keyboard/_0583_ ;
wire \keyboard/_0584_ ;
wire \keyboard/_0585_ ;
wire \keyboard/_0586_ ;
wire \keyboard/_0587_ ;
wire \keyboard/_0588_ ;
wire \keyboard/_0589_ ;
wire \keyboard/_0590_ ;
wire \keyboard/_0591_ ;
wire \keyboard/_0592_ ;
wire \keyboard/_0593_ ;
wire \keyboard/_0594_ ;
wire \keyboard/_0595_ ;
wire \keyboard/_0596_ ;
wire \keyboard/_0597_ ;
wire \keyboard/_0598_ ;
wire \keyboard/_0599_ ;
wire \keyboard/_0600_ ;
wire \keyboard/_0601_ ;
wire \keyboard/_0602_ ;
wire \keyboard/_0603_ ;
wire \keyboard/_0604_ ;
wire \keyboard/_0605_ ;
wire \keyboard/_0606_ ;
wire \keyboard/_0607_ ;
wire \keyboard/_0608_ ;
wire \keyboard/_0609_ ;
wire \keyboard/_0610_ ;
wire \keyboard/_0611_ ;
wire \keyboard/_0612_ ;
wire \keyboard/_0613_ ;
wire \keyboard/_0614_ ;
wire \keyboard/_0615_ ;
wire \keyboard/_0616_ ;
wire \keyboard/_0617_ ;
wire \keyboard/_0618_ ;
wire \keyboard/_0619_ ;
wire \keyboard/_0620_ ;
wire \keyboard/_0621_ ;
wire \keyboard/_0622_ ;
wire \keyboard/_0623_ ;
wire \keyboard/_0624_ ;
wire \keyboard/_0625_ ;
wire \keyboard/_0626_ ;
wire \keyboard/_0627_ ;
wire \keyboard/_0628_ ;
wire \keyboard/_0629_ ;
wire \keyboard/_0630_ ;
wire \keyboard/_0631_ ;
wire \keyboard/_0632_ ;
wire \keyboard/_0633_ ;
wire \keyboard/_0634_ ;
wire \keyboard/_0635_ ;
wire \keyboard/_0636_ ;
wire \keyboard/_0637_ ;
wire \keyboard/_0638_ ;
wire \keyboard/_0639_ ;
wire \keyboard/_0640_ ;
wire \keyboard/_0641_ ;
wire \keyboard/_0642_ ;
wire \keyboard/_0643_ ;
wire \keyboard/_0644_ ;
wire \keyboard/_0645_ ;
wire \keyboard/_0646_ ;
wire \keyboard/_0647_ ;
wire \keyboard/_0648_ ;
wire \keyboard/_0649_ ;
wire \keyboard/_0650_ ;
wire \keyboard/_0651_ ;
wire \keyboard/_0652_ ;
wire \keyboard/_0653_ ;
wire \keyboard/_0654_ ;
wire \keyboard/_0655_ ;
wire \keyboard/_0656_ ;
wire \keyboard/_0657_ ;
wire \keyboard/_0658_ ;
wire \keyboard/_0659_ ;
wire \keyboard/_0660_ ;
wire \keyboard/_0661_ ;
wire \keyboard/_0662_ ;
wire \keyboard/_0663_ ;
wire \keyboard/_0664_ ;
wire \keyboard/_0665_ ;
wire \keyboard/_0666_ ;
wire \keyboard/_0667_ ;
wire \keyboard/_0668_ ;
wire \keyboard/_0669_ ;
wire \keyboard/_0670_ ;
wire \keyboard/_0671_ ;
wire \keyboard/_0672_ ;
wire \keyboard/_0673_ ;
wire \keyboard/_0674_ ;
wire \keyboard/_0675_ ;
wire \keyboard/_0676_ ;
wire \keyboard/_0677_ ;
wire \keyboard/_0678_ ;
wire \keyboard/_0679_ ;
wire \keyboard/_0680_ ;
wire \keyboard/_0681_ ;
wire \keyboard/_0682_ ;
wire \keyboard/_0683_ ;
wire \keyboard/_0684_ ;
wire \keyboard/_0685_ ;
wire \keyboard/_0686_ ;
wire \keyboard/_0687_ ;
wire \keyboard/_0688_ ;
wire \keyboard/_0689_ ;
wire \keyboard/_0690_ ;
wire \keyboard/_0691_ ;
wire \keyboard/_0692_ ;
wire \keyboard/_0693_ ;
wire \keyboard/_0694_ ;
wire \keyboard/_0695_ ;
wire \keyboard/_0696_ ;
wire \keyboard/_0697_ ;
wire \keyboard/_0698_ ;
wire \keyboard/_0699_ ;
wire \keyboard/_0700_ ;
wire \keyboard/_0701_ ;
wire \keyboard/_0702_ ;
wire \keyboard/_0703_ ;
wire \keyboard/_0704_ ;
wire \keyboard/_0705_ ;
wire \keyboard/_0706_ ;
wire \keyboard/_0707_ ;
wire \keyboard/_0708_ ;
wire \keyboard/_0709_ ;
wire \keyboard/_0710_ ;
wire \keyboard/_0711_ ;
wire \keyboard/_0712_ ;
wire \keyboard/_0713_ ;
wire \keyboard/_0714_ ;
wire \keyboard/_0715_ ;
wire \keyboard/_0716_ ;
wire \keyboard/_0717_ ;
wire \keyboard/_0718_ ;
wire \keyboard/_0719_ ;
wire \keyboard/_0720_ ;
wire \keyboard/_0721_ ;
wire \keyboard/_0722_ ;
wire \keyboard/_0723_ ;
wire \keyboard/_0724_ ;
wire \keyboard/_0725_ ;
wire \keyboard/_0726_ ;
wire \keyboard/_0727_ ;
wire \keyboard/_0728_ ;
wire \keyboard/_0729_ ;
wire \keyboard/_0730_ ;
wire \keyboard/_0731_ ;
wire \keyboard/_0732_ ;
wire \keyboard/_0733_ ;
wire \keyboard/_0734_ ;
wire \keyboard/_0735_ ;
wire \keyboard/_0736_ ;
wire \keyboard/_0737_ ;
wire \keyboard/_0738_ ;
wire \keyboard/_0739_ ;
wire \keyboard/_0740_ ;
wire \keyboard/_0741_ ;
wire \keyboard/_0742_ ;
wire \keyboard/_0743_ ;
wire \keyboard/_0744_ ;
wire \keyboard/_0745_ ;
wire \keyboard/_0746_ ;
wire \keyboard/_0747_ ;
wire \keyboard/_0748_ ;
wire \keyboard/_0749_ ;
wire \keyboard/_0750_ ;
wire \keyboard/_0751_ ;
wire \keyboard/_0752_ ;
wire \keyboard/_0753_ ;
wire \keyboard/_0754_ ;
wire \keyboard/_0755_ ;
wire \keyboard/_0756_ ;
wire \keyboard/_0757_ ;
wire \keyboard/_0758_ ;
wire \keyboard/_0759_ ;
wire \keyboard/_0760_ ;
wire \keyboard/_0761_ ;
wire \keyboard/_0762_ ;
wire \keyboard/_0763_ ;
wire \seg0/_000_ ;
wire \seg0/_001_ ;
wire \seg0/_002_ ;
wire \seg0/_003_ ;
wire \seg0/_004_ ;
wire \seg0/_005_ ;
wire \seg0/_006_ ;
wire \seg0/_007_ ;
wire \seg0/_008_ ;
wire \seg0/_009_ ;
wire \seg0/_010_ ;
wire \seg0/_011_ ;
wire \seg0/_012_ ;
wire \seg0/_013_ ;
wire \seg0/_014_ ;
wire \seg0/_015_ ;
wire \seg0/_016_ ;
wire \seg0/_017_ ;
wire \seg0/_018_ ;
wire \seg0/_019_ ;
wire \seg0/_020_ ;
wire \seg0/_021_ ;
wire \seg0/_022_ ;
wire \seg0/_023_ ;
wire \seg0/_024_ ;
wire \seg0/_025_ ;
wire \seg0/_026_ ;
wire \seg0/_027_ ;
wire \seg0/_028_ ;
wire \seg0/_029_ ;
wire \seg0/_030_ ;
wire \seg0/_031_ ;
wire \seg0/_032_ ;
wire \seg0/_033_ ;
wire \seg0/_034_ ;
wire \seg0/_035_ ;
wire \seg0/_036_ ;
wire \seg0/_037_ ;
wire \seg0/_038_ ;
wire \seg0/_039_ ;
wire \seg0/_040_ ;
wire \seg0/_041_ ;
wire \seg0/_042_ ;
wire \seg0/_043_ ;
wire \seg0/_044_ ;
wire \seg0/_045_ ;
wire \seg0/_046_ ;
wire \seg0/_047_ ;
wire \seg0/_048_ ;
wire \seg0/_049_ ;
wire \seg0/_050_ ;
wire \seg0/_051_ ;
wire \seg0/_052_ ;
wire \seg0/_053_ ;
wire \seg0/_054_ ;
wire \seg0/_055_ ;
wire \seg0/_056_ ;
wire \seg0/_057_ ;
wire \seg0/_058_ ;
wire \seg0/_059_ ;
wire \seg0/_060_ ;
wire \seg0/_061_ ;
wire \seg1/_000_ ;
wire \seg1/_001_ ;
wire \seg1/_002_ ;
wire \seg1/_003_ ;
wire \seg1/_004_ ;
wire \seg1/_005_ ;
wire \seg1/_006_ ;
wire \seg1/_007_ ;
wire \seg1/_008_ ;
wire \seg1/_009_ ;
wire \seg1/_010_ ;
wire \seg1/_011_ ;
wire \seg1/_012_ ;
wire \seg1/_013_ ;
wire \seg1/_014_ ;
wire \seg1/_015_ ;
wire \seg1/_016_ ;
wire \seg1/_017_ ;
wire \seg1/_018_ ;
wire \seg1/_019_ ;
wire \seg1/_020_ ;
wire \seg1/_021_ ;
wire \seg1/_022_ ;
wire \seg1/_023_ ;
wire \seg1/_024_ ;
wire \seg1/_025_ ;
wire \seg1/_026_ ;
wire \seg1/_027_ ;
wire \seg1/_028_ ;
wire \seg1/_029_ ;
wire \seg1/_030_ ;
wire \seg1/_031_ ;
wire \seg1/_032_ ;
wire \seg1/_033_ ;
wire \seg1/_034_ ;
wire \seg1/_035_ ;
wire \seg1/_036_ ;
wire \seg1/_037_ ;
wire \seg1/_038_ ;
wire \seg1/_039_ ;
wire \seg1/_040_ ;
wire \seg1/_041_ ;
wire \seg1/_042_ ;
wire \seg1/_043_ ;
wire \seg1/_044_ ;
wire \seg1/_045_ ;
wire \seg1/_046_ ;
wire \seg1/_047_ ;
wire \seg1/_048_ ;
wire \seg1/_049_ ;
wire \seg1/_050_ ;
wire \seg1/_051_ ;
wire \seg1/_052_ ;
wire \seg1/_053_ ;
wire \seg1/_054_ ;
wire \seg1/_055_ ;
wire \seg1/_056_ ;
wire \seg1/_057_ ;
wire \seg1/_058_ ;
wire \seg1/_059_ ;
wire \seg1/_060_ ;
wire \seg1/_061_ ;
wire \seg2/_000_ ;
wire \seg2/_001_ ;
wire \seg2/_002_ ;
wire \seg2/_003_ ;
wire \seg2/_004_ ;
wire \seg2/_005_ ;
wire \seg2/_006_ ;
wire \seg2/_007_ ;
wire \seg2/_008_ ;
wire \seg2/_009_ ;
wire \seg2/_010_ ;
wire \seg2/_011_ ;
wire \seg2/_012_ ;
wire \seg2/_013_ ;
wire \seg2/_014_ ;
wire \seg2/_015_ ;
wire \seg2/_016_ ;
wire \seg2/_017_ ;
wire \seg2/_018_ ;
wire \seg2/_019_ ;
wire \seg2/_020_ ;
wire \seg2/_021_ ;
wire \seg2/_022_ ;
wire \seg2/_023_ ;
wire \seg2/_024_ ;
wire \seg2/_025_ ;
wire \seg2/_026_ ;
wire \seg2/_027_ ;
wire \seg2/_028_ ;
wire \seg2/_029_ ;
wire \seg2/_030_ ;
wire \seg2/_031_ ;
wire \seg2/_032_ ;
wire \seg2/_033_ ;
wire \seg2/_034_ ;
wire \seg2/_035_ ;
wire \seg2/_036_ ;
wire \seg2/_037_ ;
wire \seg2/_038_ ;
wire \seg2/_039_ ;
wire \seg2/_040_ ;
wire \seg2/_041_ ;
wire \seg2/_042_ ;
wire \seg2/_043_ ;
wire \seg2/_044_ ;
wire \seg2/_045_ ;
wire \seg2/_046_ ;
wire \seg2/_047_ ;
wire \seg2/_048_ ;
wire \seg2/_049_ ;
wire \seg2/_050_ ;
wire \seg2/_051_ ;
wire \seg2/_052_ ;
wire \seg2/_053_ ;
wire \seg2/_054_ ;
wire \seg2/_055_ ;
wire \seg2/_056_ ;
wire \seg2/_057_ ;
wire \seg2/_058_ ;
wire \seg2/_059_ ;
wire \seg2/_060_ ;
wire \seg2/_061_ ;
wire \seg3/_000_ ;
wire \seg3/_001_ ;
wire \seg3/_002_ ;
wire \seg3/_003_ ;
wire \seg3/_004_ ;
wire \seg3/_005_ ;
wire \seg3/_006_ ;
wire \seg3/_007_ ;
wire \seg3/_008_ ;
wire \seg3/_009_ ;
wire \seg3/_010_ ;
wire \seg3/_011_ ;
wire \seg3/_012_ ;
wire \seg3/_013_ ;
wire \seg3/_014_ ;
wire \seg3/_015_ ;
wire \seg3/_016_ ;
wire \seg3/_017_ ;
wire \seg3/_018_ ;
wire \seg3/_019_ ;
wire \seg3/_020_ ;
wire \seg3/_021_ ;
wire \seg3/_022_ ;
wire \seg3/_023_ ;
wire \seg3/_024_ ;
wire \seg3/_025_ ;
wire \seg3/_026_ ;
wire \seg3/_027_ ;
wire \seg3/_028_ ;
wire \seg3/_029_ ;
wire \seg3/_030_ ;
wire \seg3/_031_ ;
wire \seg3/_032_ ;
wire \seg3/_033_ ;
wire \seg3/_034_ ;
wire \seg3/_035_ ;
wire \seg3/_036_ ;
wire \seg3/_037_ ;
wire \seg3/_038_ ;
wire \seg3/_039_ ;
wire \seg3/_040_ ;
wire \seg3/_041_ ;
wire \seg3/_042_ ;
wire \seg3/_043_ ;
wire \seg3/_044_ ;
wire \seg3/_045_ ;
wire \seg3/_046_ ;
wire \seg3/_047_ ;
wire \seg3/_048_ ;
wire \seg3/_049_ ;
wire \seg3/_050_ ;
wire \seg3/_051_ ;
wire \seg3/_052_ ;
wire \seg3/_053_ ;
wire \seg3/_054_ ;
wire \seg3/_055_ ;
wire \seg3/_056_ ;
wire \seg3/_057_ ;
wire \seg3/_058_ ;
wire \seg3/_059_ ;
wire \seg3/_060_ ;
wire \seg3/_061_ ;
wire \seg4/_000_ ;
wire \seg4/_001_ ;
wire \seg4/_002_ ;
wire \seg4/_003_ ;
wire \seg4/_004_ ;
wire \seg4/_005_ ;
wire \seg4/_006_ ;
wire \seg4/_007_ ;
wire \seg4/_008_ ;
wire \seg4/_009_ ;
wire \seg4/_010_ ;
wire \seg4/_011_ ;
wire \seg4/_012_ ;
wire \seg4/_013_ ;
wire \seg4/_014_ ;
wire \seg4/_015_ ;
wire \seg4/_016_ ;
wire \seg4/_017_ ;
wire \seg4/_018_ ;
wire \seg4/_019_ ;
wire \seg4/_020_ ;
wire \seg4/_021_ ;
wire \seg4/_022_ ;
wire \seg4/_023_ ;
wire \seg4/_024_ ;
wire \seg4/_025_ ;
wire \seg4/_026_ ;
wire \seg4/_027_ ;
wire \seg4/_028_ ;
wire \seg4/_029_ ;
wire \seg4/_030_ ;
wire \seg4/_031_ ;
wire \seg4/_032_ ;
wire \seg4/_033_ ;
wire \seg4/_034_ ;
wire \seg4/_035_ ;
wire \seg4/_036_ ;
wire \seg4/_037_ ;
wire \seg4/_038_ ;
wire \seg4/_039_ ;
wire \seg4/_040_ ;
wire \seg4/_041_ ;
wire \seg4/_042_ ;
wire \seg4/_043_ ;
wire \seg4/_044_ ;
wire \seg4/_045_ ;
wire \seg4/_046_ ;
wire \seg4/_047_ ;
wire \seg4/_048_ ;
wire \seg4/_049_ ;
wire \seg4/_050_ ;
wire \seg4/_051_ ;
wire \seg4/_052_ ;
wire \seg4/_053_ ;
wire \seg4/_054_ ;
wire \seg4/_055_ ;
wire \seg4/_056_ ;
wire \seg4/_057_ ;
wire \seg4/_058_ ;
wire \seg4/_059_ ;
wire \seg4/_060_ ;
wire \seg4/_061_ ;
wire \seg5/_000_ ;
wire \seg5/_001_ ;
wire \seg5/_002_ ;
wire \seg5/_003_ ;
wire \seg5/_004_ ;
wire \seg5/_005_ ;
wire \seg5/_006_ ;
wire \seg5/_007_ ;
wire \seg5/_008_ ;
wire \seg5/_009_ ;
wire \seg5/_010_ ;
wire \seg5/_011_ ;
wire \seg5/_012_ ;
wire \seg5/_013_ ;
wire \seg5/_014_ ;
wire \seg5/_015_ ;
wire \seg5/_016_ ;
wire \seg5/_017_ ;
wire \seg5/_018_ ;
wire \seg5/_019_ ;
wire \seg5/_020_ ;
wire \seg5/_021_ ;
wire \seg5/_022_ ;
wire \seg5/_023_ ;
wire \seg5/_024_ ;
wire \seg5/_025_ ;
wire \seg5/_026_ ;
wire \seg5/_027_ ;
wire \seg5/_028_ ;
wire \seg5/_029_ ;
wire \seg5/_030_ ;
wire \seg5/_031_ ;
wire \seg5/_032_ ;
wire \seg5/_033_ ;
wire \seg5/_034_ ;
wire \seg5/_035_ ;
wire \seg5/_036_ ;
wire \seg5/_037_ ;
wire \seg5/_038_ ;
wire \seg5/_039_ ;
wire \seg5/_040_ ;
wire \seg5/_041_ ;
wire \seg5/_042_ ;
wire \seg5/_043_ ;
wire \seg5/_044_ ;
wire \seg5/_045_ ;
wire \seg5/_046_ ;
wire \seg5/_047_ ;
wire \seg5/_048_ ;
wire \seg5/_049_ ;
wire \seg5/_050_ ;
wire \seg5/_051_ ;
wire \seg5/_052_ ;
wire \seg5/_053_ ;
wire \seg5/_054_ ;
wire \seg5/_055_ ;
wire \seg5/_056_ ;
wire \seg5/_057_ ;
wire \seg5/_058_ ;
wire \seg5/_059_ ;
wire \seg5/_060_ ;
wire \seg5/_061_ ;
wire reset ;
wire io_clrn ;
wire clock ;
wire io_ps2_clk ;
wire io_ps2_data ;
wire \counter_io_ones[0] ;
wire \counter_io_ones[1] ;
wire \counter_io_ones[2] ;
wire \counter_io_ones[3] ;
wire \counter_io_tens[0] ;
wire \counter_io_tens[1] ;
wire \counter_io_tens[2] ;
wire \counter_io_tens[3] ;
wire \data_d1[0] ;
wire \data_d1[1] ;
wire \data_d1[2] ;
wire \data_d1[3] ;
wire \data_d1[4] ;
wire \data_d1[5] ;
wire \data_d1[6] ;
wire \data_d1[7] ;
wire \decoder_io_ascii[0] ;
wire \decoder_io_ascii[1] ;
wire \decoder_io_ascii[2] ;
wire \decoder_io_ascii[3] ;
wire \decoder_io_ascii[4] ;
wire \decoder_io_ascii[5] ;
wire \decoder_io_ascii[6] ;
wire \decoder_io_ascii[7] ;
wire \key_ascii_display_reg[0] ;
wire \key_ascii_display_reg[1] ;
wire \key_ascii_display_reg[2] ;
wire \key_ascii_display_reg[3] ;
wire \key_ascii_display_reg[4] ;
wire \key_ascii_display_reg[5] ;
wire \key_ascii_display_reg[6] ;
wire \key_ascii_display_reg[7] ;
wire \key_scan_display_reg[0] ;
wire \key_scan_display_reg[1] ;
wire \key_scan_display_reg[2] ;
wire \key_scan_display_reg[3] ;
wire \key_scan_display_reg[4] ;
wire \key_scan_display_reg[5] ;
wire \key_scan_display_reg[6] ;
wire \key_scan_display_reg[7] ;
wire \keyboard_io_data[0] ;
wire \keyboard_io_data[1] ;
wire \keyboard_io_data[2] ;
wire \keyboard_io_data[3] ;
wire \keyboard_io_data[4] ;
wire \keyboard_io_data[5] ;
wire \keyboard_io_data[6] ;
wire \keyboard_io_data[7] ;
wire \seg0_in[0] ;
wire \seg0_in[1] ;
wire \seg0_in[2] ;
wire \seg0_in[3] ;
wire \seg1_in[0] ;
wire \seg1_in[1] ;
wire \seg1_in[2] ;
wire \seg1_in[3] ;
wire \seg2_in[0] ;
wire \seg2_in[1] ;
wire \seg2_in[2] ;
wire \seg2_in[3] ;
wire \seg3_in[0] ;
wire \seg3_in[1] ;
wire \seg3_in[2] ;
wire \seg3_in[3] ;
wire \keyboard/_ps2_clk_sync_T_1[0] ;
wire \keyboard/_ps2_clk_sync_T_1[1] ;
wire \keyboard/_ps2_clk_sync_T_1[2] ;
wire \keyboard/buffer[0] ;
wire \keyboard/buffer[1] ;
wire \keyboard/buffer[2] ;
wire \keyboard/buffer[3] ;
wire \keyboard/buffer[4] ;
wire \keyboard/buffer[5] ;
wire \keyboard/buffer[6] ;
wire \keyboard/buffer[7] ;
wire \keyboard/buffer[8] ;
wire \keyboard/buffer[9] ;
wire \keyboard/count[0] ;
wire \keyboard/count[1] ;
wire \keyboard/count[2] ;
wire \keyboard/count[3] ;
wire \keyboard/fifo_0[0] ;
wire \keyboard/fifo_0[1] ;
wire \keyboard/fifo_0[2] ;
wire \keyboard/fifo_0[3] ;
wire \keyboard/fifo_0[4] ;
wire \keyboard/fifo_0[5] ;
wire \keyboard/fifo_0[6] ;
wire \keyboard/fifo_0[7] ;
wire \keyboard/fifo_1[0] ;
wire \keyboard/fifo_1[1] ;
wire \keyboard/fifo_1[2] ;
wire \keyboard/fifo_1[3] ;
wire \keyboard/fifo_1[4] ;
wire \keyboard/fifo_1[5] ;
wire \keyboard/fifo_1[6] ;
wire \keyboard/fifo_1[7] ;
wire \keyboard/fifo_2[0] ;
wire \keyboard/fifo_2[1] ;
wire \keyboard/fifo_2[2] ;
wire \keyboard/fifo_2[3] ;
wire \keyboard/fifo_2[4] ;
wire \keyboard/fifo_2[5] ;
wire \keyboard/fifo_2[6] ;
wire \keyboard/fifo_2[7] ;
wire \keyboard/fifo_3[0] ;
wire \keyboard/fifo_3[1] ;
wire \keyboard/fifo_3[2] ;
wire \keyboard/fifo_3[3] ;
wire \keyboard/fifo_3[4] ;
wire \keyboard/fifo_3[5] ;
wire \keyboard/fifo_3[6] ;
wire \keyboard/fifo_3[7] ;
wire \keyboard/fifo_4[0] ;
wire \keyboard/fifo_4[1] ;
wire \keyboard/fifo_4[2] ;
wire \keyboard/fifo_4[3] ;
wire \keyboard/fifo_4[4] ;
wire \keyboard/fifo_4[5] ;
wire \keyboard/fifo_4[6] ;
wire \keyboard/fifo_4[7] ;
wire \keyboard/fifo_5[0] ;
wire \keyboard/fifo_5[1] ;
wire \keyboard/fifo_5[2] ;
wire \keyboard/fifo_5[3] ;
wire \keyboard/fifo_5[4] ;
wire \keyboard/fifo_5[5] ;
wire \keyboard/fifo_5[6] ;
wire \keyboard/fifo_5[7] ;
wire \keyboard/fifo_6[0] ;
wire \keyboard/fifo_6[1] ;
wire \keyboard/fifo_6[2] ;
wire \keyboard/fifo_6[3] ;
wire \keyboard/fifo_6[4] ;
wire \keyboard/fifo_6[5] ;
wire \keyboard/fifo_6[6] ;
wire \keyboard/fifo_6[7] ;
wire \keyboard/fifo_7[0] ;
wire \keyboard/fifo_7[1] ;
wire \keyboard/fifo_7[2] ;
wire \keyboard/fifo_7[3] ;
wire \keyboard/fifo_7[4] ;
wire \keyboard/fifo_7[5] ;
wire \keyboard/fifo_7[6] ;
wire \keyboard/fifo_7[7] ;
wire \keyboard/ps2_clk_sync[0] ;
wire \keyboard/ps2_clk_sync[1] ;
wire \keyboard/ps2_clk_sync[2] ;
wire \keyboard/r_ptr[0] ;
wire \keyboard/r_ptr[1] ;
wire \keyboard/r_ptr[2] ;
wire \keyboard/w_ptr[0] ;
wire \keyboard/w_ptr[1] ;
wire \keyboard/w_ptr[2] ;
wire \io_seg_out_0[0] ;
wire \io_seg_out_0[1] ;
wire \io_seg_out_0[2] ;
wire \io_seg_out_0[3] ;
wire \io_seg_out_0[4] ;
wire \io_seg_out_0[5] ;
wire \io_seg_out_0[6] ;
wire \io_seg_out_0[7] ;
wire \io_seg_out_1[0] ;
wire \io_seg_out_1[1] ;
wire \io_seg_out_1[2] ;
wire \io_seg_out_1[3] ;
wire \io_seg_out_1[4] ;
wire \io_seg_out_1[5] ;
wire \io_seg_out_1[6] ;
wire \io_seg_out_1[7] ;
wire \io_seg_out_2[0] ;
wire \io_seg_out_2[1] ;
wire \io_seg_out_2[2] ;
wire \io_seg_out_2[3] ;
wire \io_seg_out_2[4] ;
wire \io_seg_out_2[5] ;
wire \io_seg_out_2[6] ;
wire \io_seg_out_2[7] ;
wire \io_seg_out_3[0] ;
wire \io_seg_out_3[1] ;
wire \io_seg_out_3[2] ;
wire \io_seg_out_3[3] ;
wire \io_seg_out_3[4] ;
wire \io_seg_out_3[5] ;
wire \io_seg_out_3[6] ;
wire \io_seg_out_3[7] ;
wire \io_seg_out_4[0] ;
wire \io_seg_out_4[1] ;
wire \io_seg_out_4[2] ;
wire \io_seg_out_4[3] ;
wire \io_seg_out_4[4] ;
wire \io_seg_out_4[5] ;
wire \io_seg_out_4[6] ;
wire \io_seg_out_4[7] ;
wire \io_seg_out_5[0] ;
wire \io_seg_out_5[1] ;
wire \io_seg_out_5[2] ;
wire \io_seg_out_5[3] ;
wire \io_seg_out_5[4] ;
wire \io_seg_out_5[5] ;
wire \io_seg_out_5[6] ;
wire \io_seg_out_5[7] ;

assign io_seg_out_0[0] = \io_seg_out_0[0] ;
assign io_seg_out_0[1] = \io_seg_out_0[1] ;
assign io_seg_out_0[2] = \io_seg_out_0[2] ;
assign io_seg_out_0[3] = \io_seg_out_0[3] ;
assign io_seg_out_0[4] = \io_seg_out_0[4] ;
assign io_seg_out_0[5] = \io_seg_out_0[5] ;
assign io_seg_out_0[6] = \io_seg_out_0[6] ;
assign io_seg_out_0[7] = \io_seg_out_0[7] ;
assign io_seg_out_1[0] = \io_seg_out_1[0] ;
assign io_seg_out_1[1] = \io_seg_out_1[1] ;
assign io_seg_out_1[2] = \io_seg_out_1[2] ;
assign io_seg_out_1[3] = \io_seg_out_1[3] ;
assign io_seg_out_1[4] = \io_seg_out_1[4] ;
assign io_seg_out_1[5] = \io_seg_out_1[5] ;
assign io_seg_out_1[6] = \io_seg_out_1[6] ;
assign io_seg_out_1[7] = \io_seg_out_1[7] ;
assign io_seg_out_2[0] = \io_seg_out_2[0] ;
assign io_seg_out_2[1] = \io_seg_out_2[1] ;
assign io_seg_out_2[2] = \io_seg_out_2[2] ;
assign io_seg_out_2[3] = \io_seg_out_2[3] ;
assign io_seg_out_2[4] = \io_seg_out_2[4] ;
assign io_seg_out_2[5] = \io_seg_out_2[5] ;
assign io_seg_out_2[6] = \io_seg_out_2[6] ;
assign io_seg_out_2[7] = \io_seg_out_2[7] ;
assign io_seg_out_3[0] = \io_seg_out_3[0] ;
assign io_seg_out_3[1] = \io_seg_out_3[1] ;
assign io_seg_out_3[2] = \io_seg_out_3[2] ;
assign io_seg_out_3[3] = \io_seg_out_3[3] ;
assign io_seg_out_3[4] = \io_seg_out_3[4] ;
assign io_seg_out_3[5] = \io_seg_out_3[5] ;
assign io_seg_out_3[6] = \io_seg_out_3[6] ;
assign io_seg_out_3[7] = \io_seg_out_3[7] ;
assign io_seg_out_4[0] = \io_seg_out_4[0] ;
assign io_seg_out_4[1] = \io_seg_out_4[1] ;
assign io_seg_out_4[2] = \io_seg_out_4[2] ;
assign io_seg_out_4[3] = \io_seg_out_4[3] ;
assign io_seg_out_4[4] = \io_seg_out_4[4] ;
assign io_seg_out_4[5] = \io_seg_out_4[5] ;
assign io_seg_out_4[6] = \io_seg_out_4[6] ;
assign io_seg_out_4[7] = \io_seg_out_4[7] ;
assign io_seg_out_5[0] = \io_seg_out_5[0] ;
assign io_seg_out_5[1] = \io_seg_out_5[1] ;
assign io_seg_out_5[2] = \io_seg_out_5[2] ;
assign io_seg_out_5[3] = \io_seg_out_5[3] ;
assign io_seg_out_5[4] = \io_seg_out_5[4] ;
assign io_seg_out_5[5] = \io_seg_out_5[5] ;
assign io_seg_out_5[6] = \io_seg_out_5[6] ;
assign io_seg_out_5[7] = \io_seg_out_5[7] ;

AND2_X1 _195_ ( .A1(_082_ ), .A2(_072_ ), .ZN(_150_ ) );
AND2_X1 _196_ ( .A1(_072_ ), .A2(_083_ ), .ZN(_151_ ) );
AND2_X1 _197_ ( .A1(_072_ ), .A2(_084_ ), .ZN(_152_ ) );
AND2_X1 _198_ ( .A1(_072_ ), .A2(_085_ ), .ZN(_153_ ) );
AND2_X1 _199_ ( .A1(_072_ ), .A2(_086_ ), .ZN(_154_ ) );
AND2_X1 _200_ ( .A1(_072_ ), .A2(_087_ ), .ZN(_155_ ) );
AND2_X1 _201_ ( .A1(_072_ ), .A2(_088_ ), .ZN(_156_ ) );
AND2_X1 _202_ ( .A1(_072_ ), .A2(_089_ ), .ZN(_157_ ) );
AND2_X1 _203_ ( .A1(_072_ ), .A2(_074_ ), .ZN(_158_ ) );
AND2_X1 _204_ ( .A1(_072_ ), .A2(_075_ ), .ZN(_159_ ) );
AND2_X1 _205_ ( .A1(_072_ ), .A2(_076_ ), .ZN(_160_ ) );
AND2_X1 _206_ ( .A1(_072_ ), .A2(_077_ ), .ZN(_161_ ) );
AND2_X1 _207_ ( .A1(_072_ ), .A2(_078_ ), .ZN(_162_ ) );
AND2_X1 _208_ ( .A1(_072_ ), .A2(_079_ ), .ZN(_163_ ) );
AND2_X1 _209_ ( .A1(_072_ ), .A2(_080_ ), .ZN(_164_ ) );
AND2_X1 _210_ ( .A1(_072_ ), .A2(_081_ ), .ZN(_165_ ) );
INV_X32 _211_ ( .A(_098_ ), .ZN(_099_ ) );
NOR2_X4 _212_ ( .A1(_099_ ), .A2(_148_ ), .ZN(_100_ ) );
BUF_X8 _213_ ( .A(_100_ ), .Z(_101_ ) );
INV_X1 _214_ ( .A(_055_ ), .ZN(_102_ ) );
AOI21_X1 _215_ ( .A(_101_ ), .B1(_072_ ), .B2(_102_ ), .ZN(_103_ ) );
INV_X1 _216_ ( .A(_149_ ), .ZN(_104_ ) );
NAND2_X2 _217_ ( .A1(_104_ ), .A2(_073_ ), .ZN(_105_ ) );
NOR2_X1 _218_ ( .A1(_103_ ), .A2(_105_ ), .ZN(_035_ ) );
MUX2_X1 _219_ ( .A(_074_ ), .B(_064_ ), .S(_101_ ), .Z(_106_ ) );
AND3_X1 _220_ ( .A1(_106_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_036_ ) );
MUX2_X1 _221_ ( .A(_075_ ), .B(_065_ ), .S(_100_ ), .Z(_107_ ) );
AND3_X1 _222_ ( .A1(_107_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_037_ ) );
MUX2_X1 _223_ ( .A(_076_ ), .B(_066_ ), .S(_100_ ), .Z(_108_ ) );
AND3_X1 _224_ ( .A1(_108_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_038_ ) );
MUX2_X1 _225_ ( .A(_077_ ), .B(_067_ ), .S(_100_ ), .Z(_109_ ) );
AND3_X1 _226_ ( .A1(_109_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_039_ ) );
MUX2_X1 _227_ ( .A(_078_ ), .B(_068_ ), .S(_100_ ), .Z(_110_ ) );
AND3_X1 _228_ ( .A1(_110_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_040_ ) );
MUX2_X1 _229_ ( .A(_079_ ), .B(_069_ ), .S(_100_ ), .Z(_111_ ) );
AND3_X1 _230_ ( .A1(_111_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_041_ ) );
MUX2_X1 _231_ ( .A(_080_ ), .B(_070_ ), .S(_100_ ), .Z(_112_ ) );
AND3_X1 _232_ ( .A1(_112_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_042_ ) );
MUX2_X1 _233_ ( .A(_081_ ), .B(_071_ ), .S(_100_ ), .Z(_113_ ) );
AND3_X1 _234_ ( .A1(_113_ ), .A2(_104_ ), .A3(_073_ ), .ZN(_043_ ) );
AND2_X1 _235_ ( .A1(_101_ ), .A2(_090_ ), .ZN(_114_ ) );
INV_X1 _236_ ( .A(_114_ ), .ZN(_115_ ) );
BUF_X4 _237_ ( .A(_099_ ), .Z(_116_ ) );
BUF_X4 _238_ ( .A(_116_ ), .Z(_117_ ) );
OAI21_X1 _239_ ( .A(_082_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_118_ ) );
AOI21_X1 _240_ ( .A(_105_ ), .B1(_115_ ), .B2(_118_ ), .ZN(_044_ ) );
AND2_X1 _241_ ( .A1(_101_ ), .A2(_091_ ), .ZN(_119_ ) );
INV_X1 _242_ ( .A(_119_ ), .ZN(_120_ ) );
OAI21_X1 _243_ ( .A(_083_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_121_ ) );
AOI21_X1 _244_ ( .A(_105_ ), .B1(_120_ ), .B2(_121_ ), .ZN(_045_ ) );
AND2_X1 _245_ ( .A1(_101_ ), .A2(_092_ ), .ZN(_122_ ) );
INV_X1 _246_ ( .A(_122_ ), .ZN(_123_ ) );
OAI21_X1 _247_ ( .A(_084_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_124_ ) );
AOI21_X1 _248_ ( .A(_105_ ), .B1(_123_ ), .B2(_124_ ), .ZN(_046_ ) );
AND2_X1 _249_ ( .A1(_101_ ), .A2(_093_ ), .ZN(_125_ ) );
INV_X1 _250_ ( .A(_125_ ), .ZN(_126_ ) );
OAI21_X1 _251_ ( .A(_085_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_127_ ) );
AOI21_X1 _252_ ( .A(_105_ ), .B1(_126_ ), .B2(_127_ ), .ZN(_047_ ) );
AND2_X1 _253_ ( .A1(_101_ ), .A2(_094_ ), .ZN(_128_ ) );
INV_X1 _254_ ( .A(_128_ ), .ZN(_129_ ) );
OAI21_X1 _255_ ( .A(_086_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_130_ ) );
AOI21_X1 _256_ ( .A(_105_ ), .B1(_129_ ), .B2(_130_ ), .ZN(_048_ ) );
AND2_X1 _257_ ( .A1(_101_ ), .A2(_095_ ), .ZN(_131_ ) );
INV_X1 _258_ ( .A(_131_ ), .ZN(_132_ ) );
OAI21_X1 _259_ ( .A(_087_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_133_ ) );
AOI21_X1 _260_ ( .A(_105_ ), .B1(_132_ ), .B2(_133_ ), .ZN(_049_ ) );
AND2_X1 _261_ ( .A1(_101_ ), .A2(_096_ ), .ZN(_134_ ) );
INV_X1 _262_ ( .A(_134_ ), .ZN(_135_ ) );
OAI21_X1 _263_ ( .A(_088_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_136_ ) );
AOI21_X1 _264_ ( .A(_105_ ), .B1(_135_ ), .B2(_136_ ), .ZN(_050_ ) );
AND2_X1 _265_ ( .A1(_101_ ), .A2(_097_ ), .ZN(_137_ ) );
INV_X1 _266_ ( .A(_137_ ), .ZN(_138_ ) );
OAI21_X1 _267_ ( .A(_089_ ), .B1(_117_ ), .B2(_148_ ), .ZN(_139_ ) );
AOI21_X1 _268_ ( .A(_105_ ), .B1(_138_ ), .B2(_139_ ), .ZN(_051_ ) );
NOR2_X1 _269_ ( .A1(_117_ ), .A2(_149_ ), .ZN(_053_ ) );
OAI21_X1 _270_ ( .A(_056_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_140_ ) );
AOI21_X1 _271_ ( .A(_149_ ), .B1(_115_ ), .B2(_140_ ), .ZN(_027_ ) );
OAI21_X1 _272_ ( .A(_057_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_141_ ) );
AOI21_X1 _273_ ( .A(_149_ ), .B1(_120_ ), .B2(_141_ ), .ZN(_028_ ) );
OAI21_X1 _274_ ( .A(_058_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_142_ ) );
AOI21_X1 _275_ ( .A(_149_ ), .B1(_123_ ), .B2(_142_ ), .ZN(_029_ ) );
OAI21_X1 _276_ ( .A(_059_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_143_ ) );
AOI21_X1 _277_ ( .A(_149_ ), .B1(_126_ ), .B2(_143_ ), .ZN(_030_ ) );
OAI21_X1 _278_ ( .A(_060_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_144_ ) );
AOI21_X1 _279_ ( .A(_149_ ), .B1(_129_ ), .B2(_144_ ), .ZN(_031_ ) );
OAI21_X1 _280_ ( .A(_061_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_145_ ) );
AOI21_X1 _281_ ( .A(_149_ ), .B1(_132_ ), .B2(_145_ ), .ZN(_032_ ) );
OAI21_X1 _282_ ( .A(_062_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_146_ ) );
AOI21_X1 _283_ ( .A(_149_ ), .B1(_135_ ), .B2(_146_ ), .ZN(_033_ ) );
OAI21_X1 _284_ ( .A(_063_ ), .B1(_116_ ), .B2(_148_ ), .ZN(_147_ ) );
AOI21_X1 _285_ ( .A(_149_ ), .B1(_138_ ), .B2(_147_ ), .ZN(_034_ ) );
NOR3_X1 _286_ ( .A1(_117_ ), .A2(_148_ ), .A3(_055_ ), .ZN(_054_ ) );
OR3_X1 _287_ ( .A1(_116_ ), .A2(_149_ ), .A3(_148_ ), .ZN(_052_ ) );
LOGIC1_X1 _288_ ( .Z(_193_ ) );
LOGIC0_X1 _289_ ( .Z(_194_ ) );
BUF_X1 _290_ ( .A(\key_scan_display_reg[0] ), .Z(_082_ ) );
BUF_X1 _291_ ( .A(display_en ), .Z(_072_ ) );
BUF_X1 _292_ ( .A(_150_ ), .Z(\seg0_in[0] ) );
BUF_X1 _293_ ( .A(\key_scan_display_reg[1] ), .Z(_083_ ) );
BUF_X1 _294_ ( .A(_151_ ), .Z(\seg0_in[1] ) );
BUF_X1 _295_ ( .A(\key_scan_display_reg[2] ), .Z(_084_ ) );
BUF_X1 _296_ ( .A(_152_ ), .Z(\seg0_in[2] ) );
BUF_X1 _297_ ( .A(\key_scan_display_reg[3] ), .Z(_085_ ) );
BUF_X1 _298_ ( .A(_153_ ), .Z(\seg0_in[3] ) );
BUF_X1 _299_ ( .A(\key_scan_display_reg[4] ), .Z(_086_ ) );
BUF_X1 _300_ ( .A(_154_ ), .Z(\seg1_in[0] ) );
BUF_X1 _301_ ( .A(\key_scan_display_reg[5] ), .Z(_087_ ) );
BUF_X1 _302_ ( .A(_155_ ), .Z(\seg1_in[1] ) );
BUF_X1 _303_ ( .A(\key_scan_display_reg[6] ), .Z(_088_ ) );
BUF_X1 _304_ ( .A(_156_ ), .Z(\seg1_in[2] ) );
BUF_X1 _305_ ( .A(\key_scan_display_reg[7] ), .Z(_089_ ) );
BUF_X1 _306_ ( .A(_157_ ), .Z(\seg1_in[3] ) );
BUF_X1 _307_ ( .A(\key_ascii_display_reg[0] ), .Z(_074_ ) );
BUF_X1 _308_ ( .A(_158_ ), .Z(\seg2_in[0] ) );
BUF_X1 _309_ ( .A(\key_ascii_display_reg[1] ), .Z(_075_ ) );
BUF_X1 _310_ ( .A(_159_ ), .Z(\seg2_in[1] ) );
BUF_X1 _311_ ( .A(\key_ascii_display_reg[2] ), .Z(_076_ ) );
BUF_X1 _312_ ( .A(_160_ ), .Z(\seg2_in[2] ) );
BUF_X1 _313_ ( .A(\key_ascii_display_reg[3] ), .Z(_077_ ) );
BUF_X1 _314_ ( .A(_161_ ), .Z(\seg2_in[3] ) );
BUF_X1 _315_ ( .A(\key_ascii_display_reg[4] ), .Z(_078_ ) );
BUF_X1 _316_ ( .A(_162_ ), .Z(\seg3_in[0] ) );
BUF_X1 _317_ ( .A(\key_ascii_display_reg[5] ), .Z(_079_ ) );
BUF_X1 _318_ ( .A(_163_ ), .Z(\seg3_in[1] ) );
BUF_X1 _319_ ( .A(\key_ascii_display_reg[6] ), .Z(_080_ ) );
BUF_X1 _320_ ( .A(_164_ ), .Z(\seg3_in[2] ) );
BUF_X1 _321_ ( .A(\key_ascii_display_reg[7] ), .Z(_081_ ) );
BUF_X1 _322_ ( .A(_165_ ), .Z(\seg3_in[3] ) );
BUF_X1 _323_ ( .A(reset ), .Z(_149_ ) );
BUF_X1 _324_ ( .A(keyboard_io_ready ), .Z(_098_ ) );
BUF_X1 _325_ ( .A(ready_delay ), .Z(_148_ ) );
BUF_X1 _326_ ( .A(counter_io_key_release ), .Z(_055_ ) );
BUF_X1 _327_ ( .A(io_clrn ), .Z(_073_ ) );
BUF_X1 _328_ ( .A(_035_ ), .Z(_008_ ) );
BUF_X1 _329_ ( .A(\decoder_io_ascii[0] ), .Z(_064_ ) );
BUF_X1 _330_ ( .A(_036_ ), .Z(_009_ ) );
BUF_X1 _331_ ( .A(\decoder_io_ascii[1] ), .Z(_065_ ) );
BUF_X1 _332_ ( .A(_037_ ), .Z(_010_ ) );
BUF_X1 _333_ ( .A(\decoder_io_ascii[2] ), .Z(_066_ ) );
BUF_X1 _334_ ( .A(_038_ ), .Z(_011_ ) );
BUF_X1 _335_ ( .A(\decoder_io_ascii[3] ), .Z(_067_ ) );
BUF_X1 _336_ ( .A(_039_ ), .Z(_012_ ) );
BUF_X1 _337_ ( .A(\decoder_io_ascii[4] ), .Z(_068_ ) );
BUF_X1 _338_ ( .A(_040_ ), .Z(_013_ ) );
BUF_X1 _339_ ( .A(\decoder_io_ascii[5] ), .Z(_069_ ) );
BUF_X1 _340_ ( .A(_041_ ), .Z(_014_ ) );
BUF_X1 _341_ ( .A(\decoder_io_ascii[6] ), .Z(_070_ ) );
BUF_X1 _342_ ( .A(_042_ ), .Z(_015_ ) );
BUF_X1 _343_ ( .A(\decoder_io_ascii[7] ), .Z(_071_ ) );
BUF_X1 _344_ ( .A(_043_ ), .Z(_016_ ) );
BUF_X1 _345_ ( .A(\keyboard_io_data[0] ), .Z(_090_ ) );
BUF_X1 _346_ ( .A(_044_ ), .Z(_017_ ) );
BUF_X1 _347_ ( .A(\keyboard_io_data[1] ), .Z(_091_ ) );
BUF_X1 _348_ ( .A(_045_ ), .Z(_018_ ) );
BUF_X1 _349_ ( .A(\keyboard_io_data[2] ), .Z(_092_ ) );
BUF_X1 _350_ ( .A(_046_ ), .Z(_019_ ) );
BUF_X1 _351_ ( .A(\keyboard_io_data[3] ), .Z(_093_ ) );
BUF_X1 _352_ ( .A(_047_ ), .Z(_020_ ) );
BUF_X1 _353_ ( .A(\keyboard_io_data[4] ), .Z(_094_ ) );
BUF_X1 _354_ ( .A(_048_ ), .Z(_021_ ) );
BUF_X1 _355_ ( .A(\keyboard_io_data[5] ), .Z(_095_ ) );
BUF_X1 _356_ ( .A(_049_ ), .Z(_022_ ) );
BUF_X1 _357_ ( .A(\keyboard_io_data[6] ), .Z(_096_ ) );
BUF_X1 _358_ ( .A(_050_ ), .Z(_023_ ) );
BUF_X1 _359_ ( .A(\keyboard_io_data[7] ), .Z(_097_ ) );
BUF_X1 _360_ ( .A(_051_ ), .Z(_024_ ) );
BUF_X1 _361_ ( .A(_053_ ), .Z(_026_ ) );
BUF_X1 _362_ ( .A(\data_d1[0] ), .Z(_056_ ) );
BUF_X1 _363_ ( .A(_027_ ), .Z(_000_ ) );
BUF_X1 _364_ ( .A(\data_d1[1] ), .Z(_057_ ) );
BUF_X1 _365_ ( .A(_028_ ), .Z(_001_ ) );
BUF_X1 _366_ ( .A(\data_d1[2] ), .Z(_058_ ) );
BUF_X1 _367_ ( .A(_029_ ), .Z(_002_ ) );
BUF_X1 _368_ ( .A(\data_d1[3] ), .Z(_059_ ) );
BUF_X1 _369_ ( .A(_030_ ), .Z(_003_ ) );
BUF_X1 _370_ ( .A(\data_d1[4] ), .Z(_060_ ) );
BUF_X1 _371_ ( .A(_031_ ), .Z(_004_ ) );
BUF_X1 _372_ ( .A(\data_d1[5] ), .Z(_061_ ) );
BUF_X1 _373_ ( .A(_032_ ), .Z(_005_ ) );
BUF_X1 _374_ ( .A(\data_d1[6] ), .Z(_062_ ) );
BUF_X1 _375_ ( .A(_033_ ), .Z(_006_ ) );
BUF_X1 _376_ ( .A(\data_d1[7] ), .Z(_063_ ) );
BUF_X1 _377_ ( .A(_034_ ), .Z(_007_ ) );
BUF_X1 _378_ ( .A(_054_ ), .Z(counter_io_key_press ) );
BUF_X1 _379_ ( .A(_052_ ), .Z(_025_ ) );
DFF_X1 _380_ ( .D(_025_ ), .CK(clock ), .Q(keyboard_io_nextdata_n ), .QN(_166_ ) );
DFF_X1 _381_ ( .D(_026_ ), .CK(clock ), .Q(ready_delay ), .QN(_167_ ) );
DFF_X1 _382_ ( .D(_000_ ), .CK(clock ), .Q(\data_d1[0] ), .QN(_168_ ) );
DFF_X1 _383_ ( .D(_001_ ), .CK(clock ), .Q(\data_d1[1] ), .QN(_169_ ) );
DFF_X1 _384_ ( .D(_002_ ), .CK(clock ), .Q(\data_d1[2] ), .QN(_170_ ) );
DFF_X1 _385_ ( .D(_003_ ), .CK(clock ), .Q(\data_d1[3] ), .QN(_171_ ) );
DFF_X1 _386_ ( .D(_004_ ), .CK(clock ), .Q(\data_d1[4] ), .QN(_172_ ) );
DFF_X1 _387_ ( .D(_005_ ), .CK(clock ), .Q(\data_d1[5] ), .QN(_173_ ) );
DFF_X1 _388_ ( .D(_006_ ), .CK(clock ), .Q(\data_d1[6] ), .QN(_174_ ) );
DFF_X1 _389_ ( .D(_007_ ), .CK(clock ), .Q(\data_d1[7] ), .QN(_175_ ) );
DFF_X1 _390_ ( .D(_017_ ), .CK(clock ), .Q(\key_scan_display_reg[0] ), .QN(_176_ ) );
DFF_X1 _391_ ( .D(_018_ ), .CK(clock ), .Q(\key_scan_display_reg[1] ), .QN(_177_ ) );
DFF_X1 _392_ ( .D(_019_ ), .CK(clock ), .Q(\key_scan_display_reg[2] ), .QN(_178_ ) );
DFF_X1 _393_ ( .D(_020_ ), .CK(clock ), .Q(\key_scan_display_reg[3] ), .QN(_179_ ) );
DFF_X1 _394_ ( .D(_021_ ), .CK(clock ), .Q(\key_scan_display_reg[4] ), .QN(_180_ ) );
DFF_X1 _395_ ( .D(_022_ ), .CK(clock ), .Q(\key_scan_display_reg[5] ), .QN(_181_ ) );
DFF_X1 _396_ ( .D(_023_ ), .CK(clock ), .Q(\key_scan_display_reg[6] ), .QN(_182_ ) );
DFF_X1 _397_ ( .D(_024_ ), .CK(clock ), .Q(\key_scan_display_reg[7] ), .QN(_183_ ) );
DFF_X1 _398_ ( .D(_009_ ), .CK(clock ), .Q(\key_ascii_display_reg[0] ), .QN(_184_ ) );
DFF_X1 _399_ ( .D(_010_ ), .CK(clock ), .Q(\key_ascii_display_reg[1] ), .QN(_185_ ) );
DFF_X1 _400_ ( .D(_011_ ), .CK(clock ), .Q(\key_ascii_display_reg[2] ), .QN(_186_ ) );
DFF_X1 _401_ ( .D(_012_ ), .CK(clock ), .Q(\key_ascii_display_reg[3] ), .QN(_187_ ) );
DFF_X1 _402_ ( .D(_013_ ), .CK(clock ), .Q(\key_ascii_display_reg[4] ), .QN(_188_ ) );
DFF_X1 _403_ ( .D(_014_ ), .CK(clock ), .Q(\key_ascii_display_reg[5] ), .QN(_189_ ) );
DFF_X1 _404_ ( .D(_015_ ), .CK(clock ), .Q(\key_ascii_display_reg[6] ), .QN(_190_ ) );
DFF_X1 _405_ ( .D(_016_ ), .CK(clock ), .Q(\key_ascii_display_reg[7] ), .QN(_191_ ) );
DFF_X1 _406_ ( .D(_008_ ), .CK(clock ), .Q(display_en ), .QN(_192_ ) );
INV_X32 \counter/_084_ ( .A(\counter/_033_ ), .ZN(\counter/_044_ ) );
NOR2_X4 \counter/_085_ ( .A1(\counter/_044_ ), .A2(\counter/_081_ ), .ZN(\counter/_045_ ) );
OAI21_X1 \counter/_086_ ( .A(\counter/_045_ ), .B1(\counter/_034_ ), .B2(\counter/_032_ ), .ZN(\counter/_046_ ) );
NOR2_X1 \counter/_087_ ( .A1(\counter/_046_ ), .A2(\counter/_035_ ), .ZN(\counter/_016_ ) );
INV_X8 \counter/_088_ ( .A(\counter/_045_ ), .ZN(\counter/_047_ ) );
INV_X16 \counter/_089_ ( .A(\counter/_036_ ), .ZN(\counter/_048_ ) );
NOR2_X4 \counter/_090_ ( .A1(\counter/_048_ ), .A2(\counter/_037_ ), .ZN(\counter/_049_ ) );
INV_X32 \counter/_091_ ( .A(\counter/_039_ ), .ZN(\counter/_050_ ) );
NOR2_X4 \counter/_092_ ( .A1(\counter/_050_ ), .A2(\counter/_038_ ), .ZN(\counter/_051_ ) );
INV_X32 \counter/_093_ ( .A(\counter/_034_ ), .ZN(\counter/_052_ ) );
NOR2_X4 \counter/_094_ ( .A1(\counter/_052_ ), .A2(\counter/_032_ ), .ZN(\counter/_053_ ) );
AND4_X1 \counter/_095_ ( .A1(\counter/_040_ ), .A2(\counter/_049_ ), .A3(\counter/_051_ ), .A4(\counter/_053_ ), .ZN(\counter/_054_ ) );
AND2_X4 \counter/_096_ ( .A1(\counter/_049_ ), .A2(\counter/_051_ ), .ZN(\counter/_055_ ) );
AND2_X4 \counter/_097_ ( .A1(\counter/_055_ ), .A2(\counter/_053_ ), .ZN(\counter/_056_ ) );
INV_X4 \counter/_098_ ( .A(\counter/_056_ ), .ZN(\counter/_057_ ) );
AOI211_X2 \counter/_099_ ( .A(\counter/_047_ ), .B(\counter/_054_ ), .C1(\counter/_057_ ), .C2(\counter/_025_ ), .ZN(\counter/_021_ ) );
INV_X1 \counter/_100_ ( .A(\counter/_041_ ), .ZN(\counter/_058_ ) );
AND3_X1 \counter/_101_ ( .A1(\counter/_058_ ), .A2(\counter/_040_ ), .A3(\counter/_043_ ), .ZN(\counter/_059_ ) );
INV_X1 \counter/_102_ ( .A(\counter/_042_ ), .ZN(\counter/_060_ ) );
NAND2_X1 \counter/_103_ ( .A1(\counter/_059_ ), .A2(\counter/_060_ ), .ZN(\counter/_061_ ) );
XOR2_X1 \counter/_104_ ( .A(\counter/_040_ ), .B(\counter/_041_ ), .Z(\counter/_062_ ) );
NAND4_X1 \counter/_105_ ( .A1(\counter/_056_ ), .A2(\counter/_045_ ), .A3(\counter/_061_ ), .A4(\counter/_062_ ), .ZN(\counter/_063_ ) );
NOR2_X2 \counter/_106_ ( .A1(\counter/_056_ ), .A2(\counter/_047_ ), .ZN(\counter/_064_ ) );
INV_X2 \counter/_107_ ( .A(\counter/_064_ ), .ZN(\counter/_065_ ) );
OAI21_X1 \counter/_108_ ( .A(\counter/_063_ ), .B1(\counter/_065_ ), .B2(\counter/_026_ ), .ZN(\counter/_022_ ) );
NAND2_X1 \counter/_109_ ( .A1(\counter/_040_ ), .A2(\counter/_041_ ), .ZN(\counter/_066_ ) );
XNOR2_X1 \counter/_110_ ( .A(\counter/_066_ ), .B(\counter/_060_ ), .ZN(\counter/_067_ ) );
AND3_X1 \counter/_111_ ( .A1(\counter/_067_ ), .A2(\counter/_055_ ), .A3(\counter/_053_ ), .ZN(\counter/_068_ ) );
AOI211_X2 \counter/_112_ ( .A(\counter/_047_ ), .B(\counter/_068_ ), .C1(\counter/_057_ ), .C2(\counter/_027_ ), .ZN(\counter/_023_ ) );
OR3_X1 \counter/_113_ ( .A1(\counter/_066_ ), .A2(\counter/_060_ ), .A3(\counter/_028_ ), .ZN(\counter/_069_ ) );
AOI21_X4 \counter/_114_ ( .A(\counter/_057_ ), .B1(\counter/_061_ ), .B2(\counter/_069_ ), .ZN(\counter/_070_ ) );
NAND4_X4 \counter/_115_ ( .A1(\counter/_056_ ), .A2(\counter/_040_ ), .A3(\counter/_041_ ), .A4(\counter/_042_ ), .ZN(\counter/_071_ ) );
AOI211_X2 \counter/_116_ ( .A(\counter/_047_ ), .B(\counter/_070_ ), .C1(\counter/_028_ ), .C2(\counter/_071_ ), .ZN(\counter/_024_ ) );
AND2_X1 \counter/_117_ ( .A1(\counter/_053_ ), .A2(\counter/_036_ ), .ZN(\counter/_072_ ) );
INV_X1 \counter/_118_ ( .A(\counter/_053_ ), .ZN(\counter/_073_ ) );
AOI211_X2 \counter/_119_ ( .A(\counter/_047_ ), .B(\counter/_072_ ), .C1(\counter/_029_ ), .C2(\counter/_073_ ), .ZN(\counter/_017_ ) );
AND2_X1 \counter/_120_ ( .A1(\counter/_048_ ), .A2(\counter/_037_ ), .ZN(\counter/_074_ ) );
NOR3_X1 \counter/_121_ ( .A1(\counter/_073_ ), .A2(\counter/_049_ ), .A3(\counter/_074_ ), .ZN(\counter/_075_ ) );
AOI211_X2 \counter/_122_ ( .A(\counter/_075_ ), .B(\counter/_065_ ), .C1(\counter/_030_ ), .C2(\counter/_073_ ), .ZN(\counter/_018_ ) );
AND3_X4 \counter/_123_ ( .A1(\counter/_053_ ), .A2(\counter/_036_ ), .A3(\counter/_037_ ), .ZN(\counter/_076_ ) );
OAI21_X1 \counter/_124_ ( .A(\counter/_045_ ), .B1(\counter/_076_ ), .B2(\counter/_038_ ), .ZN(\counter/_077_ ) );
AOI21_X1 \counter/_125_ ( .A(\counter/_077_ ), .B1(\counter/_038_ ), .B2(\counter/_076_ ), .ZN(\counter/_019_ ) );
INV_X1 \counter/_126_ ( .A(\counter/_031_ ), .ZN(\counter/_078_ ) );
AND3_X1 \counter/_127_ ( .A1(\counter/_076_ ), .A2(\counter/_038_ ), .A3(\counter/_078_ ), .ZN(\counter/_079_ ) );
AOI21_X1 \counter/_128_ ( .A(\counter/_078_ ), .B1(\counter/_076_ ), .B2(\counter/_038_ ), .ZN(\counter/_080_ ) );
NOR4_X1 \counter/_129_ ( .A1(\counter/_079_ ), .A2(\counter/_080_ ), .A3(\counter/_056_ ), .A4(\counter/_047_ ), .ZN(\counter/_020_ ) );
BUF_X1 \counter/_130_ ( .A(reset ), .Z(\counter/_081_ ) );
BUF_X1 \counter/_131_ ( .A(io_clrn ), .Z(\counter/_033_ ) );
BUF_X1 \counter/_132_ ( .A(counter_io_key_press ), .Z(\counter/_034_ ) );
BUF_X1 \counter/_133_ ( .A(\counter/counted ), .Z(\counter/_032_ ) );
BUF_X1 \counter/_134_ ( .A(counter_io_key_release ), .Z(\counter/_035_ ) );
BUF_X1 \counter/_135_ ( .A(\counter/_016_ ), .Z(\counter/_000_ ) );
BUF_X1 \counter/_136_ ( .A(\counter_io_tens[0] ), .Z(\counter/_040_ ) );
BUF_X1 \counter/_137_ ( .A(\counter_io_tens[1] ), .Z(\counter/_041_ ) );
BUF_X1 \counter/_138_ ( .A(\counter_io_tens[3] ), .Z(\counter/_043_ ) );
BUF_X1 \counter/_139_ ( .A(\counter_io_tens[2] ), .Z(\counter/_042_ ) );
BUF_X1 \counter/_140_ ( .A(\counter_io_ones[0] ), .Z(\counter/_036_ ) );
BUF_X1 \counter/_141_ ( .A(\counter_io_ones[1] ), .Z(\counter/_037_ ) );
BUF_X1 \counter/_142_ ( .A(\counter_io_ones[3] ), .Z(\counter/_039_ ) );
BUF_X1 \counter/_143_ ( .A(\counter_io_ones[2] ), .Z(\counter/_038_ ) );
BUF_X1 \counter/_144_ ( .A(\counter/_009_ ), .Z(\counter/_025_ ) );
BUF_X1 \counter/_145_ ( .A(\counter/_021_ ), .Z(\counter/_005_ ) );
BUF_X1 \counter/_146_ ( .A(\counter/_010_ ), .Z(\counter/_026_ ) );
BUF_X1 \counter/_147_ ( .A(\counter/_022_ ), .Z(\counter/_006_ ) );
BUF_X1 \counter/_148_ ( .A(\counter/_011_ ), .Z(\counter/_027_ ) );
BUF_X1 \counter/_149_ ( .A(\counter/_023_ ), .Z(\counter/_007_ ) );
BUF_X1 \counter/_150_ ( .A(\counter/_012_ ), .Z(\counter/_028_ ) );
BUF_X1 \counter/_151_ ( .A(\counter/_024_ ), .Z(\counter/_008_ ) );
BUF_X1 \counter/_152_ ( .A(\counter/_013_ ), .Z(\counter/_029_ ) );
BUF_X1 \counter/_153_ ( .A(\counter/_017_ ), .Z(\counter/_001_ ) );
BUF_X1 \counter/_154_ ( .A(\counter/_014_ ), .Z(\counter/_030_ ) );
BUF_X1 \counter/_155_ ( .A(\counter/_018_ ), .Z(\counter/_002_ ) );
BUF_X1 \counter/_156_ ( .A(\counter/_019_ ), .Z(\counter/_003_ ) );
BUF_X1 \counter/_157_ ( .A(\counter/_015_ ), .Z(\counter/_031_ ) );
BUF_X1 \counter/_158_ ( .A(\counter/_020_ ), .Z(\counter/_004_ ) );
DFF_X1 \counter/_159_ ( .D(\counter/_001_ ), .CK(clock ), .Q(\counter_io_ones[0] ), .QN(\counter/_013_ ) );
DFF_X1 \counter/_160_ ( .D(\counter/_002_ ), .CK(clock ), .Q(\counter_io_ones[1] ), .QN(\counter/_014_ ) );
DFF_X1 \counter/_161_ ( .D(\counter/_003_ ), .CK(clock ), .Q(\counter_io_ones[2] ), .QN(\counter/_082_ ) );
DFF_X1 \counter/_162_ ( .D(\counter/_004_ ), .CK(clock ), .Q(\counter_io_ones[3] ), .QN(\counter/_015_ ) );
DFF_X1 \counter/_163_ ( .D(\counter/_005_ ), .CK(clock ), .Q(\counter_io_tens[0] ), .QN(\counter/_009_ ) );
DFF_X1 \counter/_164_ ( .D(\counter/_006_ ), .CK(clock ), .Q(\counter_io_tens[1] ), .QN(\counter/_010_ ) );
DFF_X1 \counter/_165_ ( .D(\counter/_007_ ), .CK(clock ), .Q(\counter_io_tens[2] ), .QN(\counter/_011_ ) );
DFF_X1 \counter/_166_ ( .D(\counter/_008_ ), .CK(clock ), .Q(\counter_io_tens[3] ), .QN(\counter/_012_ ) );
DFF_X1 \counter/_167_ ( .D(\counter/_000_ ), .CK(clock ), .Q(\counter/counted ), .QN(\counter/_083_ ) );
INV_X1 \decoder/_133_ ( .A(\decoder/_011_ ), .ZN(\decoder/_055_ ) );
OR2_X1 \decoder/_134_ ( .A1(\decoder/_055_ ), .A2(\decoder/_021_ ), .ZN(\decoder/_056_ ) );
INV_X32 \decoder/_135_ ( .A(\decoder/_017_ ), .ZN(\decoder/_057_ ) );
NOR2_X4 \decoder/_136_ ( .A1(\decoder/_057_ ), .A2(\decoder/_016_ ), .ZN(\decoder/_058_ ) );
NOR2_X4 \decoder/_137_ ( .A1(\decoder/_018_ ), .A2(\decoder/_019_ ), .ZN(\decoder/_059_ ) );
AND2_X4 \decoder/_138_ ( .A1(\decoder/_058_ ), .A2(\decoder/_059_ ), .ZN(\decoder/_060_ ) );
AND2_X4 \decoder/_139_ ( .A1(\decoder/_015_ ), .A2(\decoder/_014_ ), .ZN(\decoder/_061_ ) );
INV_X1 \decoder/_140_ ( .A(\decoder/_012_ ), .ZN(\decoder/_062_ ) );
AND3_X1 \decoder/_141_ ( .A1(\decoder/_061_ ), .A2(\decoder/_062_ ), .A3(\decoder/_013_ ), .ZN(\decoder/_063_ ) );
AND2_X1 \decoder/_142_ ( .A1(\decoder/_060_ ), .A2(\decoder/_063_ ), .ZN(\decoder/_064_ ) );
NOR2_X1 \decoder/_143_ ( .A1(\decoder/_062_ ), .A2(\decoder/_013_ ), .ZN(\decoder/_065_ ) );
AND2_X4 \decoder/_144_ ( .A1(\decoder/_065_ ), .A2(\decoder/_061_ ), .ZN(\decoder/_066_ ) );
AND2_X4 \decoder/_145_ ( .A1(\decoder/_017_ ), .A2(\decoder/_016_ ), .ZN(\decoder/_067_ ) );
AND2_X4 \decoder/_146_ ( .A1(\decoder/_067_ ), .A2(\decoder/_059_ ), .ZN(\decoder/_068_ ) );
AND2_X1 \decoder/_147_ ( .A1(\decoder/_066_ ), .A2(\decoder/_068_ ), .ZN(\decoder/_069_ ) );
NOR2_X1 \decoder/_148_ ( .A1(\decoder/_064_ ), .A2(\decoder/_069_ ), .ZN(\decoder/_070_ ) );
INV_X1 \decoder/_149_ ( .A(\decoder/_070_ ), .ZN(\decoder/_071_ ) );
INV_X16 \decoder/_150_ ( .A(\decoder/_015_ ), .ZN(\decoder/_072_ ) );
AND2_X4 \decoder/_151_ ( .A1(\decoder/_072_ ), .A2(\decoder/_014_ ), .ZN(\decoder/_073_ ) );
INV_X32 \decoder/_152_ ( .A(\decoder/_013_ ), .ZN(\decoder/_074_ ) );
NOR2_X1 \decoder/_153_ ( .A1(\decoder/_074_ ), .A2(\decoder/_012_ ), .ZN(\decoder/_075_ ) );
AND2_X2 \decoder/_154_ ( .A1(\decoder/_073_ ), .A2(\decoder/_075_ ), .ZN(\decoder/_076_ ) );
AND2_X2 \decoder/_155_ ( .A1(\decoder/_057_ ), .A2(\decoder/_016_ ), .ZN(\decoder/_077_ ) );
AND2_X4 \decoder/_156_ ( .A1(\decoder/_077_ ), .A2(\decoder/_059_ ), .ZN(\decoder/_078_ ) );
AND2_X1 \decoder/_157_ ( .A1(\decoder/_076_ ), .A2(\decoder/_078_ ), .ZN(\decoder/_079_ ) );
BUF_X8 \decoder/_158_ ( .A(\decoder/_060_ ), .Z(\decoder/_080_ ) );
AND2_X1 \decoder/_159_ ( .A1(\decoder/_076_ ), .A2(\decoder/_080_ ), .ZN(\decoder/_081_ ) );
NOR3_X2 \decoder/_160_ ( .A1(\decoder/_071_ ), .A2(\decoder/_079_ ), .A3(\decoder/_081_ ), .ZN(\decoder/_082_ ) );
NOR2_X1 \decoder/_161_ ( .A1(\decoder/_012_ ), .A2(\decoder/_013_ ), .ZN(\decoder/_083_ ) );
AND2_X4 \decoder/_162_ ( .A1(\decoder/_073_ ), .A2(\decoder/_083_ ), .ZN(\decoder/_084_ ) );
INV_X1 \decoder/_163_ ( .A(\decoder/_018_ ), .ZN(\decoder/_085_ ) );
NOR2_X1 \decoder/_164_ ( .A1(\decoder/_085_ ), .A2(\decoder/_019_ ), .ZN(\decoder/_086_ ) );
NOR2_X1 \decoder/_165_ ( .A1(\decoder/_017_ ), .A2(\decoder/_016_ ), .ZN(\decoder/_087_ ) );
AND2_X2 \decoder/_166_ ( .A1(\decoder/_086_ ), .A2(\decoder/_087_ ), .ZN(\decoder/_088_ ) );
AND2_X1 \decoder/_167_ ( .A1(\decoder/_084_ ), .A2(\decoder/_088_ ), .ZN(\decoder/_089_ ) );
NOR2_X1 \decoder/_168_ ( .A1(\decoder/_072_ ), .A2(\decoder/_014_ ), .ZN(\decoder/_090_ ) );
AND2_X1 \decoder/_169_ ( .A1(\decoder/_090_ ), .A2(\decoder/_075_ ), .ZN(\decoder/_091_ ) );
AND2_X1 \decoder/_170_ ( .A1(\decoder/_091_ ), .A2(\decoder/_068_ ), .ZN(\decoder/_092_ ) );
NOR2_X1 \decoder/_171_ ( .A1(\decoder/_089_ ), .A2(\decoder/_092_ ), .ZN(\decoder/_093_ ) );
NOR2_X1 \decoder/_172_ ( .A1(\decoder/_015_ ), .A2(\decoder/_014_ ), .ZN(\decoder/_094_ ) );
NAND3_X1 \decoder/_173_ ( .A1(\decoder/_088_ ), .A2(\decoder/_013_ ), .A3(\decoder/_094_ ), .ZN(\decoder/_095_ ) );
AND2_X1 \decoder/_174_ ( .A1(\decoder/_093_ ), .A2(\decoder/_095_ ), .ZN(\decoder/_096_ ) );
NOR3_X1 \decoder/_175_ ( .A1(\decoder/_057_ ), .A2(\decoder/_018_ ), .A3(\decoder/_019_ ), .ZN(\decoder/_097_ ) );
AND2_X1 \decoder/_176_ ( .A1(\decoder/_084_ ), .A2(\decoder/_097_ ), .ZN(\decoder/_098_ ) );
AND3_X1 \decoder/_177_ ( .A1(\decoder/_094_ ), .A2(\decoder/_012_ ), .A3(\decoder/_074_ ), .ZN(\decoder/_099_ ) );
AND2_X2 \decoder/_178_ ( .A1(\decoder/_080_ ), .A2(\decoder/_099_ ), .ZN(\decoder/_100_ ) );
AND2_X1 \decoder/_179_ ( .A1(\decoder/_061_ ), .A2(\decoder/_083_ ), .ZN(\decoder/_101_ ) );
AND3_X1 \decoder/_180_ ( .A1(\decoder/_101_ ), .A2(\decoder/_059_ ), .A3(\decoder/_077_ ), .ZN(\decoder/_102_ ) );
NOR3_X1 \decoder/_181_ ( .A1(\decoder/_098_ ), .A2(\decoder/_100_ ), .A3(\decoder/_102_ ), .ZN(\decoder/_103_ ) );
AND3_X1 \decoder/_182_ ( .A1(\decoder/_082_ ), .A2(\decoder/_096_ ), .A3(\decoder/_103_ ), .ZN(\decoder/_104_ ) );
AOI22_X1 \decoder/_183_ ( .A1(\decoder/_078_ ), .A2(\decoder/_066_ ), .B1(\decoder/_076_ ), .B2(\decoder/_088_ ), .ZN(\decoder/_105_ ) );
AND2_X1 \decoder/_184_ ( .A1(\decoder/_073_ ), .A2(\decoder/_065_ ), .ZN(\decoder/_106_ ) );
AND2_X1 \decoder/_185_ ( .A1(\decoder/_012_ ), .A2(\decoder/_013_ ), .ZN(\decoder/_107_ ) );
AND2_X2 \decoder/_186_ ( .A1(\decoder/_090_ ), .A2(\decoder/_107_ ), .ZN(\decoder/_108_ ) );
OAI21_X1 \decoder/_187_ ( .A(\decoder/_078_ ), .B1(\decoder/_106_ ), .B2(\decoder/_108_ ), .ZN(\decoder/_109_ ) );
AND2_X2 \decoder/_188_ ( .A1(\decoder/_075_ ), .A2(\decoder/_094_ ), .ZN(\decoder/_110_ ) );
BUF_X8 \decoder/_189_ ( .A(\decoder/_068_ ), .Z(\decoder/_111_ ) );
AOI22_X1 \decoder/_190_ ( .A1(\decoder/_080_ ), .A2(\decoder/_110_ ), .B1(\decoder/_111_ ), .B2(\decoder/_101_ ), .ZN(\decoder/_112_ ) );
AND3_X1 \decoder/_191_ ( .A1(\decoder/_105_ ), .A2(\decoder/_109_ ), .A3(\decoder/_112_ ), .ZN(\decoder/_113_ ) );
AOI21_X1 \decoder/_192_ ( .A(\decoder/_056_ ), .B1(\decoder/_104_ ), .B2(\decoder/_113_ ), .ZN(\decoder/_004_ ) );
NAND2_X1 \decoder/_193_ ( .A1(\decoder/_078_ ), .A2(\decoder/_108_ ), .ZN(\decoder/_114_ ) );
AND2_X1 \decoder/_194_ ( .A1(\decoder/_066_ ), .A2(\decoder/_060_ ), .ZN(\decoder/_115_ ) );
AOI221_X1 \decoder/_195_ ( .A(\decoder/_115_ ), .B1(\decoder/_078_ ), .B2(\decoder/_084_ ), .C1(\decoder/_111_ ), .C2(\decoder/_099_ ), .ZN(\decoder/_116_ ) );
NAND2_X1 \decoder/_196_ ( .A1(\decoder/_078_ ), .A2(\decoder/_063_ ), .ZN(\decoder/_117_ ) );
AOI22_X1 \decoder/_197_ ( .A1(\decoder/_076_ ), .A2(\decoder/_111_ ), .B1(\decoder/_108_ ), .B2(\decoder/_097_ ), .ZN(\decoder/_118_ ) );
AND4_X1 \decoder/_198_ ( .A1(\decoder/_114_ ), .A2(\decoder/_116_ ), .A3(\decoder/_117_ ), .A4(\decoder/_118_ ), .ZN(\decoder/_119_ ) );
AND2_X1 \decoder/_199_ ( .A1(\decoder/_078_ ), .A2(\decoder/_066_ ), .ZN(\decoder/_120_ ) );
AND2_X1 \decoder/_200_ ( .A1(\decoder/_091_ ), .A2(\decoder/_060_ ), .ZN(\decoder/_121_ ) );
NOR2_X1 \decoder/_201_ ( .A1(\decoder/_120_ ), .A2(\decoder/_121_ ), .ZN(\decoder/_122_ ) );
AOI221_X1 \decoder/_202_ ( .A(\decoder/_069_ ), .B1(\decoder/_076_ ), .B2(\decoder/_080_ ), .C1(\decoder/_111_ ), .C2(\decoder/_110_ ), .ZN(\decoder/_123_ ) );
AOI22_X1 \decoder/_203_ ( .A1(\decoder/_084_ ), .A2(\decoder/_111_ ), .B1(\decoder/_080_ ), .B2(\decoder/_099_ ), .ZN(\decoder/_124_ ) );
OAI21_X1 \decoder/_204_ ( .A(\decoder/_088_ ), .B1(\decoder/_084_ ), .B2(\decoder/_110_ ), .ZN(\decoder/_125_ ) );
AND4_X1 \decoder/_205_ ( .A1(\decoder/_122_ ), .A2(\decoder/_123_ ), .A3(\decoder/_124_ ), .A4(\decoder/_125_ ), .ZN(\decoder/_126_ ) );
AOI21_X1 \decoder/_206_ ( .A(\decoder/_056_ ), .B1(\decoder/_119_ ), .B2(\decoder/_126_ ), .ZN(\decoder/_005_ ) );
OAI211_X2 \decoder/_207_ ( .A(\decoder/_101_ ), .B(\decoder/_059_ ), .C1(\decoder/_067_ ), .C2(\decoder/_058_ ), .ZN(\decoder/_127_ ) );
NAND2_X1 \decoder/_208_ ( .A1(\decoder/_122_ ), .A2(\decoder/_127_ ), .ZN(\decoder/_128_ ) );
AND2_X1 \decoder/_209_ ( .A1(\decoder/_108_ ), .A2(\decoder/_080_ ), .ZN(\decoder/_129_ ) );
AND2_X1 \decoder/_210_ ( .A1(\decoder/_106_ ), .A2(\decoder/_080_ ), .ZN(\decoder/_130_ ) );
AND2_X1 \decoder/_211_ ( .A1(\decoder/_107_ ), .A2(\decoder/_094_ ), .ZN(\decoder/_022_ ) );
AND2_X1 \decoder/_212_ ( .A1(\decoder/_080_ ), .A2(\decoder/_022_ ), .ZN(\decoder/_023_ ) );
NOR4_X1 \decoder/_213_ ( .A1(\decoder/_128_ ), .A2(\decoder/_129_ ), .A3(\decoder/_130_ ), .A4(\decoder/_023_ ), .ZN(\decoder/_024_ ) );
AOI22_X1 \decoder/_214_ ( .A1(\decoder/_076_ ), .A2(\decoder/_111_ ), .B1(\decoder/_084_ ), .B2(\decoder/_097_ ), .ZN(\decoder/_025_ ) );
AOI22_X1 \decoder/_215_ ( .A1(\decoder/_108_ ), .A2(\decoder/_088_ ), .B1(\decoder/_099_ ), .B2(\decoder/_111_ ), .ZN(\decoder/_026_ ) );
AND4_X1 \decoder/_216_ ( .A1(\decoder/_093_ ), .A2(\decoder/_070_ ), .A3(\decoder/_025_ ), .A4(\decoder/_026_ ), .ZN(\decoder/_027_ ) );
AOI21_X1 \decoder/_217_ ( .A(\decoder/_056_ ), .B1(\decoder/_024_ ), .B2(\decoder/_027_ ), .ZN(\decoder/_006_ ) );
OAI21_X1 \decoder/_218_ ( .A(\decoder/_111_ ), .B1(\decoder/_108_ ), .B2(\decoder/_099_ ), .ZN(\decoder/_028_ ) );
AOI22_X1 \decoder/_219_ ( .A1(\decoder/_108_ ), .A2(\decoder/_088_ ), .B1(\decoder/_111_ ), .B2(\decoder/_022_ ), .ZN(\decoder/_029_ ) );
NAND3_X1 \decoder/_220_ ( .A1(\decoder/_096_ ), .A2(\decoder/_028_ ), .A3(\decoder/_029_ ), .ZN(\decoder/_030_ ) );
AOI22_X1 \decoder/_221_ ( .A1(\decoder/_078_ ), .A2(\decoder/_084_ ), .B1(\decoder/_060_ ), .B2(\decoder/_110_ ), .ZN(\decoder/_031_ ) );
NAND3_X1 \decoder/_222_ ( .A1(\decoder/_091_ ), .A2(\decoder/_059_ ), .A3(\decoder/_077_ ), .ZN(\decoder/_032_ ) );
NAND2_X1 \decoder/_223_ ( .A1(\decoder/_031_ ), .A2(\decoder/_032_ ), .ZN(\decoder/_033_ ) );
NAND2_X1 \decoder/_224_ ( .A1(\decoder/_076_ ), .A2(\decoder/_088_ ), .ZN(\decoder/_034_ ) );
NAND2_X1 \decoder/_225_ ( .A1(\decoder/_063_ ), .A2(\decoder/_068_ ), .ZN(\decoder/_035_ ) );
NAND2_X1 \decoder/_226_ ( .A1(\decoder/_034_ ), .A2(\decoder/_035_ ), .ZN(\decoder/_036_ ) );
NOR3_X1 \decoder/_227_ ( .A1(\decoder/_030_ ), .A2(\decoder/_033_ ), .A3(\decoder/_036_ ), .ZN(\decoder/_037_ ) );
NOR2_X1 \decoder/_228_ ( .A1(\decoder/_037_ ), .A2(\decoder/_056_ ), .ZN(\decoder/_007_ ) );
INV_X1 \decoder/_229_ ( .A(\decoder/_003_ ), .ZN(\decoder/_038_ ) );
OAI21_X1 \decoder/_230_ ( .A(\decoder/_106_ ), .B1(\decoder/_088_ ), .B2(\decoder/_080_ ), .ZN(\decoder/_039_ ) );
NAND2_X1 \decoder/_231_ ( .A1(\decoder/_076_ ), .A2(\decoder/_068_ ), .ZN(\decoder/_040_ ) );
NAND3_X1 \decoder/_232_ ( .A1(\decoder/_039_ ), .A2(\decoder/_040_ ), .A3(\decoder/_117_ ), .ZN(\decoder/_041_ ) );
NOR2_X1 \decoder/_233_ ( .A1(\decoder/_041_ ), .A2(\decoder/_036_ ), .ZN(\decoder/_042_ ) );
AOI211_X2 \decoder/_234_ ( .A(\decoder/_055_ ), .B(\decoder/_038_ ), .C1(\decoder/_082_ ), .C2(\decoder/_042_ ), .ZN(\decoder/_009_ ) );
NOR2_X2 \decoder/_235_ ( .A1(\decoder/_128_ ), .A2(\decoder/_033_ ), .ZN(\decoder/_043_ ) );
OAI21_X1 \decoder/_236_ ( .A(\decoder/_066_ ), .B1(\decoder/_088_ ), .B2(\decoder/_080_ ), .ZN(\decoder/_044_ ) );
AND2_X1 \decoder/_237_ ( .A1(\decoder/_109_ ), .A2(\decoder/_044_ ), .ZN(\decoder/_045_ ) );
AOI211_X2 \decoder/_238_ ( .A(\decoder/_055_ ), .B(\decoder/_038_ ), .C1(\decoder/_043_ ), .C2(\decoder/_045_ ), .ZN(\decoder/_046_ ) );
OR2_X1 \decoder/_239_ ( .A1(\decoder/_009_ ), .A2(\decoder/_046_ ), .ZN(\decoder/_008_ ) );
INV_X1 \decoder/_240_ ( .A(\decoder/_103_ ), .ZN(\decoder/_047_ ) );
AND2_X4 \decoder/_241_ ( .A1(\decoder/_110_ ), .A2(\decoder/_111_ ), .ZN(\decoder/_048_ ) );
OR2_X4 \decoder/_242_ ( .A1(\decoder/_129_ ), .A2(\decoder/_048_ ), .ZN(\decoder/_049_ ) );
NOR4_X2 \decoder/_243_ ( .A1(\decoder/_030_ ), .A2(\decoder/_047_ ), .A3(\decoder/_023_ ), .A4(\decoder/_049_ ), .ZN(\decoder/_050_ ) );
AND2_X1 \decoder/_244_ ( .A1(\decoder/_043_ ), .A2(\decoder/_045_ ), .ZN(\decoder/_051_ ) );
AOI21_X1 \decoder/_245_ ( .A(\decoder/_056_ ), .B1(\decoder/_050_ ), .B2(\decoder/_051_ ), .ZN(\decoder/_010_ ) );
AND4_X1 \decoder/_246_ ( .A1(\decoder/_018_ ), .A2(\decoder/_019_ ), .A3(\decoder/_017_ ), .A4(\decoder/_016_ ), .ZN(\decoder/_052_ ) );
AND3_X1 \decoder/_247_ ( .A1(\decoder/_052_ ), .A2(\decoder/_083_ ), .A3(\decoder/_094_ ), .ZN(\decoder/_053_ ) );
INV_X1 \decoder/_248_ ( .A(\decoder/_053_ ), .ZN(\decoder/_054_ ) );
NOR3_X1 \decoder/_249_ ( .A1(\decoder/_054_ ), .A2(\decoder/_055_ ), .A3(\decoder/_131_ ), .ZN(\decoder/_002_ ) );
NOR3_X1 \decoder/_250_ ( .A1(\decoder/_053_ ), .A2(\decoder/_055_ ), .A3(\decoder/_003_ ), .ZN(\decoder/_020_ ) );
LOGIC0_X1 \decoder/_251_ ( .Z(\decoder/_132_ ) );
BUF_X1 \decoder/_252_ ( .A(\decoder/_132_ ), .Z(\decoder_io_ascii[7] ) );
BUF_X1 \decoder/_253_ ( .A(\data_d1[6] ), .Z(\decoder/_018_ ) );
BUF_X1 \decoder/_254_ ( .A(\data_d1[7] ), .Z(\decoder/_019_ ) );
BUF_X1 \decoder/_255_ ( .A(\data_d1[5] ), .Z(\decoder/_017_ ) );
BUF_X1 \decoder/_256_ ( .A(\data_d1[4] ), .Z(\decoder/_016_ ) );
BUF_X1 \decoder/_257_ ( .A(\data_d1[0] ), .Z(\decoder/_012_ ) );
BUF_X1 \decoder/_258_ ( .A(\data_d1[1] ), .Z(\decoder/_013_ ) );
BUF_X1 \decoder/_259_ ( .A(\data_d1[3] ), .Z(\decoder/_015_ ) );
BUF_X1 \decoder/_260_ ( .A(\data_d1[2] ), .Z(\decoder/_014_ ) );
BUF_X1 \decoder/_261_ ( .A(\decoder/isBreakCode ), .Z(\decoder/_021_ ) );
BUF_X1 \decoder/_262_ ( .A(io_clrn ), .Z(\decoder/_011_ ) );
BUF_X1 \decoder/_263_ ( .A(\decoder/_004_ ), .Z(\decoder_io_ascii[0] ) );
BUF_X1 \decoder/_264_ ( .A(\decoder/_005_ ), .Z(\decoder_io_ascii[1] ) );
BUF_X1 \decoder/_265_ ( .A(\decoder/_006_ ), .Z(\decoder_io_ascii[2] ) );
BUF_X1 \decoder/_266_ ( .A(\decoder/_007_ ), .Z(\decoder_io_ascii[3] ) );
BUF_X1 \decoder/_267_ ( .A(\decoder/_001_ ), .Z(\decoder/_003_ ) );
BUF_X1 \decoder/_268_ ( .A(\decoder/_008_ ), .Z(\decoder_io_ascii[4] ) );
BUF_X1 \decoder/_269_ ( .A(\decoder/_009_ ), .Z(\decoder_io_ascii[5] ) );
BUF_X1 \decoder/_270_ ( .A(\decoder/_010_ ), .Z(\decoder_io_ascii[6] ) );
BUF_X1 \decoder/_271_ ( .A(reset ), .Z(\decoder/_131_ ) );
BUF_X1 \decoder/_272_ ( .A(\decoder/_002_ ), .Z(\decoder/_000_ ) );
BUF_X1 \decoder/_273_ ( .A(\decoder/_020_ ), .Z(counter_io_key_release ) );
DFF_X1 \decoder/_274_ ( .D(\decoder/_000_ ), .CK(clock ), .Q(\decoder/isBreakCode ), .QN(\decoder/_001_ ) );
INV_X32 \keyboard/_0764_ ( .A(\keyboard/_0750_ ), .ZN(\keyboard/_0431_ ) );
NOR2_X4 \keyboard/_0765_ ( .A1(\keyboard/_0431_ ), .A2(\keyboard/_0751_ ), .ZN(\keyboard/_0432_ ) );
AND2_X4 \keyboard/_0766_ ( .A1(\keyboard/_0432_ ), .A2(\keyboard/_0259_ ), .ZN(\keyboard/_0433_ ) );
BUF_X8 \keyboard/_0767_ ( .A(\keyboard/_0433_ ), .Z(\keyboard/_0434_ ) );
MUX2_X1 \keyboard/_0768_ ( .A(\keyboard/_0354_ ), .B(\keyboard/_0362_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0435_ ) );
INV_X32 \keyboard/_0769_ ( .A(\keyboard/_0751_ ), .ZN(\keyboard/_0436_ ) );
NOR2_X4 \keyboard/_0770_ ( .A1(\keyboard/_0436_ ), .A2(\keyboard/_0750_ ), .ZN(\keyboard/_0437_ ) );
NAND2_X1 \keyboard/_0771_ ( .A1(\keyboard/_0437_ ), .A2(\keyboard/_0259_ ), .ZN(\keyboard/_0438_ ) );
MUX2_X2 \keyboard/_0772_ ( .A(\keyboard/_0370_ ), .B(\keyboard/_0435_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0439_ ) );
AND2_X4 \keyboard/_0773_ ( .A1(\keyboard/_0751_ ), .A2(\keyboard/_0750_ ), .ZN(\keyboard/_0440_ ) );
NAND2_X4 \keyboard/_0774_ ( .A1(\keyboard/_0440_ ), .A2(\keyboard/_0259_ ), .ZN(\keyboard/_0441_ ) );
MUX2_X2 \keyboard/_0775_ ( .A(\keyboard/_0378_ ), .B(\keyboard/_0439_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0442_ ) );
NAND2_X4 \keyboard/_0776_ ( .A1(\keyboard/_0431_ ), .A2(\keyboard/_0752_ ), .ZN(\keyboard/_0443_ ) );
NOR2_X2 \keyboard/_0777_ ( .A1(\keyboard/_0443_ ), .A2(\keyboard/_0751_ ), .ZN(\keyboard/_0444_ ) );
INV_X16 \keyboard/_0778_ ( .A(\keyboard/_0444_ ), .ZN(\keyboard/_0445_ ) );
MUX2_X2 \keyboard/_0779_ ( .A(\keyboard/_0386_ ), .B(\keyboard/_0442_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0446_ ) );
AND2_X1 \keyboard/_0780_ ( .A1(\keyboard/_0432_ ), .A2(\keyboard/_0752_ ), .ZN(\keyboard/_0447_ ) );
INV_X8 \keyboard/_0781_ ( .A(\keyboard/_0447_ ), .ZN(\keyboard/_0448_ ) );
MUX2_X2 \keyboard/_0782_ ( .A(\keyboard/_0394_ ), .B(\keyboard/_0446_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0449_ ) );
AND2_X1 \keyboard/_0783_ ( .A1(\keyboard/_0437_ ), .A2(\keyboard/_0752_ ), .ZN(\keyboard/_0450_ ) );
BUF_X32 \keyboard/_0784_ ( .A(\keyboard/_0450_ ), .Z(\keyboard/_0451_ ) );
MUX2_X2 \keyboard/_0785_ ( .A(\keyboard/_0449_ ), .B(\keyboard/_0402_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0452_ ) );
AND2_X1 \keyboard/_0786_ ( .A1(\keyboard/_0440_ ), .A2(\keyboard/_0752_ ), .ZN(\keyboard/_0453_ ) );
INV_X2 \keyboard/_0787_ ( .A(\keyboard/_0453_ ), .ZN(\keyboard/_0454_ ) );
MUX2_X2 \keyboard/_0788_ ( .A(\keyboard/_0410_ ), .B(\keyboard/_0452_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0419_ ) );
MUX2_X1 \keyboard/_0789_ ( .A(\keyboard/_0355_ ), .B(\keyboard/_0363_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0455_ ) );
MUX2_X2 \keyboard/_0790_ ( .A(\keyboard/_0371_ ), .B(\keyboard/_0455_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0456_ ) );
MUX2_X2 \keyboard/_0791_ ( .A(\keyboard/_0379_ ), .B(\keyboard/_0456_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0457_ ) );
MUX2_X2 \keyboard/_0792_ ( .A(\keyboard/_0387_ ), .B(\keyboard/_0457_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0458_ ) );
MUX2_X2 \keyboard/_0793_ ( .A(\keyboard/_0395_ ), .B(\keyboard/_0458_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0459_ ) );
MUX2_X2 \keyboard/_0794_ ( .A(\keyboard/_0459_ ), .B(\keyboard/_0403_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0460_ ) );
MUX2_X2 \keyboard/_0795_ ( .A(\keyboard/_0411_ ), .B(\keyboard/_0460_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0420_ ) );
MUX2_X1 \keyboard/_0796_ ( .A(\keyboard/_0356_ ), .B(\keyboard/_0364_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0461_ ) );
MUX2_X2 \keyboard/_0797_ ( .A(\keyboard/_0372_ ), .B(\keyboard/_0461_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0462_ ) );
MUX2_X2 \keyboard/_0798_ ( .A(\keyboard/_0380_ ), .B(\keyboard/_0462_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0463_ ) );
MUX2_X2 \keyboard/_0799_ ( .A(\keyboard/_0388_ ), .B(\keyboard/_0463_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0464_ ) );
MUX2_X2 \keyboard/_0800_ ( .A(\keyboard/_0396_ ), .B(\keyboard/_0464_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0465_ ) );
MUX2_X2 \keyboard/_0801_ ( .A(\keyboard/_0465_ ), .B(\keyboard/_0404_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0466_ ) );
MUX2_X2 \keyboard/_0802_ ( .A(\keyboard/_0412_ ), .B(\keyboard/_0466_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0421_ ) );
MUX2_X1 \keyboard/_0803_ ( .A(\keyboard/_0357_ ), .B(\keyboard/_0365_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0467_ ) );
MUX2_X2 \keyboard/_0804_ ( .A(\keyboard/_0373_ ), .B(\keyboard/_0467_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0468_ ) );
MUX2_X2 \keyboard/_0805_ ( .A(\keyboard/_0381_ ), .B(\keyboard/_0468_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0469_ ) );
MUX2_X2 \keyboard/_0806_ ( .A(\keyboard/_0389_ ), .B(\keyboard/_0469_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0470_ ) );
MUX2_X2 \keyboard/_0807_ ( .A(\keyboard/_0397_ ), .B(\keyboard/_0470_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0471_ ) );
MUX2_X2 \keyboard/_0808_ ( .A(\keyboard/_0471_ ), .B(\keyboard/_0405_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0472_ ) );
MUX2_X2 \keyboard/_0809_ ( .A(\keyboard/_0413_ ), .B(\keyboard/_0472_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0422_ ) );
MUX2_X1 \keyboard/_0810_ ( .A(\keyboard/_0358_ ), .B(\keyboard/_0366_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0473_ ) );
MUX2_X2 \keyboard/_0811_ ( .A(\keyboard/_0374_ ), .B(\keyboard/_0473_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0474_ ) );
MUX2_X2 \keyboard/_0812_ ( .A(\keyboard/_0382_ ), .B(\keyboard/_0474_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0475_ ) );
MUX2_X2 \keyboard/_0813_ ( .A(\keyboard/_0390_ ), .B(\keyboard/_0475_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0476_ ) );
MUX2_X2 \keyboard/_0814_ ( .A(\keyboard/_0398_ ), .B(\keyboard/_0476_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0477_ ) );
MUX2_X2 \keyboard/_0815_ ( .A(\keyboard/_0477_ ), .B(\keyboard/_0406_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0478_ ) );
MUX2_X2 \keyboard/_0816_ ( .A(\keyboard/_0414_ ), .B(\keyboard/_0478_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0423_ ) );
MUX2_X1 \keyboard/_0817_ ( .A(\keyboard/_0359_ ), .B(\keyboard/_0367_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0479_ ) );
MUX2_X2 \keyboard/_0818_ ( .A(\keyboard/_0375_ ), .B(\keyboard/_0479_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0480_ ) );
MUX2_X2 \keyboard/_0819_ ( .A(\keyboard/_0383_ ), .B(\keyboard/_0480_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0481_ ) );
MUX2_X2 \keyboard/_0820_ ( .A(\keyboard/_0391_ ), .B(\keyboard/_0481_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0482_ ) );
MUX2_X2 \keyboard/_0821_ ( .A(\keyboard/_0399_ ), .B(\keyboard/_0482_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0483_ ) );
MUX2_X2 \keyboard/_0822_ ( .A(\keyboard/_0483_ ), .B(\keyboard/_0407_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0484_ ) );
MUX2_X2 \keyboard/_0823_ ( .A(\keyboard/_0415_ ), .B(\keyboard/_0484_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0424_ ) );
MUX2_X1 \keyboard/_0824_ ( .A(\keyboard/_0360_ ), .B(\keyboard/_0368_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0485_ ) );
MUX2_X2 \keyboard/_0825_ ( .A(\keyboard/_0376_ ), .B(\keyboard/_0485_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0486_ ) );
MUX2_X2 \keyboard/_0826_ ( .A(\keyboard/_0384_ ), .B(\keyboard/_0486_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0487_ ) );
MUX2_X2 \keyboard/_0827_ ( .A(\keyboard/_0392_ ), .B(\keyboard/_0487_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0488_ ) );
MUX2_X2 \keyboard/_0828_ ( .A(\keyboard/_0400_ ), .B(\keyboard/_0488_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0489_ ) );
MUX2_X2 \keyboard/_0829_ ( .A(\keyboard/_0489_ ), .B(\keyboard/_0408_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0490_ ) );
MUX2_X2 \keyboard/_0830_ ( .A(\keyboard/_0416_ ), .B(\keyboard/_0490_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0425_ ) );
MUX2_X1 \keyboard/_0831_ ( .A(\keyboard/_0361_ ), .B(\keyboard/_0369_ ), .S(\keyboard/_0434_ ), .Z(\keyboard/_0491_ ) );
MUX2_X2 \keyboard/_0832_ ( .A(\keyboard/_0377_ ), .B(\keyboard/_0491_ ), .S(\keyboard/_0438_ ), .Z(\keyboard/_0492_ ) );
MUX2_X2 \keyboard/_0833_ ( .A(\keyboard/_0385_ ), .B(\keyboard/_0492_ ), .S(\keyboard/_0441_ ), .Z(\keyboard/_0493_ ) );
MUX2_X2 \keyboard/_0834_ ( .A(\keyboard/_0393_ ), .B(\keyboard/_0493_ ), .S(\keyboard/_0445_ ), .Z(\keyboard/_0494_ ) );
MUX2_X2 \keyboard/_0835_ ( .A(\keyboard/_0401_ ), .B(\keyboard/_0494_ ), .S(\keyboard/_0448_ ), .Z(\keyboard/_0495_ ) );
MUX2_X2 \keyboard/_0836_ ( .A(\keyboard/_0495_ ), .B(\keyboard/_0409_ ), .S(\keyboard/_0451_ ), .Z(\keyboard/_0496_ ) );
MUX2_X2 \keyboard/_0837_ ( .A(\keyboard/_0417_ ), .B(\keyboard/_0496_ ), .S(\keyboard/_0454_ ), .Z(\keyboard/_0426_ ) );
INV_X32 \keyboard/_0838_ ( .A(\keyboard/_0753_ ), .ZN(\keyboard/_0497_ ) );
AND2_X1 \keyboard/_0839_ ( .A1(\keyboard/_0497_ ), .A2(\keyboard/_0428_ ), .ZN(\keyboard/_0247_ ) );
AND2_X1 \keyboard/_0840_ ( .A1(\keyboard/_0497_ ), .A2(\keyboard/_0257_ ), .ZN(\keyboard/_0248_ ) );
INV_X32 \keyboard/_0841_ ( .A(\keyboard/_0258_ ), .ZN(\keyboard/_0498_ ) );
NOR2_X1 \keyboard/_0842_ ( .A1(\keyboard/_0498_ ), .A2(\keyboard/_0753_ ), .ZN(\keyboard/_0249_ ) );
AND2_X4 \keyboard/_0843_ ( .A1(\keyboard/_0497_ ), .A2(\keyboard/_0418_ ), .ZN(\keyboard/_0499_ ) );
INV_X1 \keyboard/_0844_ ( .A(\keyboard/_0499_ ), .ZN(\keyboard/_0500_ ) );
BUF_X4 \keyboard/_0845_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0501_ ) );
XOR2_X2 \keyboard/_0846_ ( .A(\keyboard/_0346_ ), .B(\keyboard/_0345_ ), .Z(\keyboard/_0502_ ) );
XNOR2_X2 \keyboard/_0847_ ( .A(\keyboard/_0344_ ), .B(\keyboard/_0343_ ), .ZN(\keyboard/_0503_ ) );
XNOR2_X2 \keyboard/_0848_ ( .A(\keyboard/_0502_ ), .B(\keyboard/_0503_ ), .ZN(\keyboard/_0504_ ) );
XOR2_X2 \keyboard/_0849_ ( .A(\keyboard/_0348_ ), .B(\keyboard/_0347_ ), .Z(\keyboard/_0505_ ) );
XNOR2_X2 \keyboard/_0850_ ( .A(\keyboard/_0342_ ), .B(\keyboard/_0341_ ), .ZN(\keyboard/_0506_ ) );
XNOR2_X2 \keyboard/_0851_ ( .A(\keyboard/_0505_ ), .B(\keyboard/_0506_ ), .ZN(\keyboard/_0507_ ) );
XNOR2_X2 \keyboard/_0852_ ( .A(\keyboard/_0504_ ), .B(\keyboard/_0507_ ), .ZN(\keyboard/_0508_ ) );
XNOR2_X2 \keyboard/_0853_ ( .A(\keyboard/_0508_ ), .B(\keyboard/_0349_ ), .ZN(\keyboard/_0509_ ) );
INV_X32 \keyboard/_0854_ ( .A(\keyboard/_0429_ ), .ZN(\keyboard/_0510_ ) );
NOR2_X1 \keyboard/_0855_ ( .A1(\keyboard/_0510_ ), .A2(\keyboard/_0340_ ), .ZN(\keyboard/_0511_ ) );
AND2_X4 \keyboard/_0856_ ( .A1(\keyboard/_0509_ ), .A2(\keyboard/_0511_ ), .ZN(\keyboard/_0512_ ) );
INV_X32 \keyboard/_0857_ ( .A(\keyboard/_0351_ ), .ZN(\keyboard/_0513_ ) );
NOR2_X4 \keyboard/_0858_ ( .A1(\keyboard/_0513_ ), .A2(\keyboard/_0350_ ), .ZN(\keyboard/_0514_ ) );
AND3_X4 \keyboard/_0859_ ( .A1(\keyboard/_0514_ ), .A2(\keyboard/_0498_ ), .A3(\keyboard/_0749_ ), .ZN(\keyboard/_0515_ ) );
INV_X16 \keyboard/_0860_ ( .A(\keyboard/_0353_ ), .ZN(\keyboard/_0516_ ) );
NOR2_X4 \keyboard/_0861_ ( .A1(\keyboard/_0516_ ), .A2(\keyboard/_0352_ ), .ZN(\keyboard/_0517_ ) );
AND2_X4 \keyboard/_0862_ ( .A1(\keyboard/_0515_ ), .A2(\keyboard/_0517_ ), .ZN(\keyboard/_0518_ ) );
NAND2_X4 \keyboard/_0863_ ( .A1(\keyboard/_0512_ ), .A2(\keyboard/_0518_ ), .ZN(\keyboard/_0519_ ) );
BUF_X16 \keyboard/_0864_ ( .A(\keyboard/_0519_ ), .Z(\keyboard/_0520_ ) );
BUF_X32 \keyboard/_0865_ ( .A(\keyboard/_0520_ ), .Z(\keyboard/_0521_ ) );
XOR2_X2 \keyboard/_0866_ ( .A(\keyboard/_0440_ ), .B(\keyboard/_0752_ ), .Z(\keyboard/_0522_ ) );
XNOR2_X1 \keyboard/_0867_ ( .A(\keyboard/_0522_ ), .B(\keyboard/_0261_ ), .ZN(\keyboard/_0523_ ) );
XNOR2_X1 \keyboard/_0868_ ( .A(\keyboard/_0751_ ), .B(\keyboard/_0750_ ), .ZN(\keyboard/_0524_ ) );
XNOR2_X1 \keyboard/_0869_ ( .A(\keyboard/_0524_ ), .B(\keyboard/_0260_ ), .ZN(\keyboard/_0525_ ) );
INV_X32 \keyboard/_0870_ ( .A(\keyboard/_0754_ ), .ZN(\keyboard/_0526_ ) );
AOI21_X1 \keyboard/_0871_ ( .A(\keyboard/_0427_ ), .B1(\keyboard/_0431_ ), .B2(\keyboard/_0526_ ), .ZN(\keyboard/_0527_ ) );
OAI211_X2 \keyboard/_0872_ ( .A(\keyboard/_0525_ ), .B(\keyboard/_0527_ ), .C1(\keyboard/_0431_ ), .C2(\keyboard/_0526_ ), .ZN(\keyboard/_0528_ ) );
OAI21_X1 \keyboard/_0873_ ( .A(\keyboard/_0430_ ), .B1(\keyboard/_0523_ ), .B2(\keyboard/_0528_ ), .ZN(\keyboard/_0529_ ) );
AOI21_X1 \keyboard/_0874_ ( .A(\keyboard/_0501_ ), .B1(\keyboard/_0521_ ), .B2(\keyboard/_0529_ ), .ZN(\keyboard/_0253_ ) );
AND2_X4 \keyboard/_0875_ ( .A1(\keyboard/_0498_ ), .A2(\keyboard/_0749_ ), .ZN(\keyboard/_0530_ ) );
AND2_X4 \keyboard/_0876_ ( .A1(\keyboard/_0530_ ), .A2(\keyboard/_0350_ ), .ZN(\keyboard/_0531_ ) );
BUF_X8 \keyboard/_0877_ ( .A(\keyboard/_0518_ ), .Z(\keyboard/_0532_ ) );
BUF_X8 \keyboard/_0878_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0533_ ) );
OR2_X4 \keyboard/_0879_ ( .A1(\keyboard/_0533_ ), .A2(\keyboard/_0500_ ), .ZN(\keyboard/_0534_ ) );
INV_X4 \keyboard/_0880_ ( .A(\keyboard/_0530_ ), .ZN(\keyboard/_0535_ ) );
AOI211_X2 \keyboard/_0881_ ( .A(\keyboard/_0531_ ), .B(\keyboard/_0534_ ), .C1(\keyboard/_0262_ ), .C2(\keyboard/_0535_ ), .ZN(\keyboard/_0179_ ) );
INV_X4 \keyboard/_0882_ ( .A(\keyboard/_0533_ ), .ZN(\keyboard/_0536_ ) );
AOI21_X2 \keyboard/_0883_ ( .A(\keyboard/_0531_ ), .B1(\keyboard/_0536_ ), .B2(\keyboard/_0351_ ), .ZN(\keyboard/_0537_ ) );
AND2_X4 \keyboard/_0884_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0351_ ), .ZN(\keyboard/_0538_ ) );
NOR3_X1 \keyboard/_0885_ ( .A1(\keyboard/_0537_ ), .A2(\keyboard/_0501_ ), .A3(\keyboard/_0538_ ), .ZN(\keyboard/_0180_ ) );
AND2_X4 \keyboard/_0886_ ( .A1(\keyboard/_0538_ ), .A2(\keyboard/_0352_ ), .ZN(\keyboard/_0539_ ) );
OAI21_X1 \keyboard/_0887_ ( .A(\keyboard/_0499_ ), .B1(\keyboard/_0538_ ), .B2(\keyboard/_0352_ ), .ZN(\keyboard/_0540_ ) );
NOR2_X1 \keyboard/_0888_ ( .A1(\keyboard/_0539_ ), .A2(\keyboard/_0540_ ), .ZN(\keyboard/_0181_ ) );
XNOR2_X2 \keyboard/_0889_ ( .A(\keyboard/_0539_ ), .B(\keyboard/_0263_ ), .ZN(\keyboard/_0541_ ) );
AND3_X1 \keyboard/_0890_ ( .A1(\keyboard/_0541_ ), .A2(\keyboard/_0536_ ), .A3(\keyboard/_0499_ ), .ZN(\keyboard/_0182_ ) );
INV_X16 \keyboard/_0891_ ( .A(\keyboard/_0427_ ), .ZN(\keyboard/_0542_ ) );
AND2_X1 \keyboard/_0892_ ( .A1(\keyboard/_0542_ ), .A2(\keyboard/_0430_ ), .ZN(\keyboard/_0543_ ) );
INV_X1 \keyboard/_0893_ ( .A(\keyboard/_0543_ ), .ZN(\keyboard/_0544_ ) );
OAI21_X1 \keyboard/_0894_ ( .A(\keyboard/_0499_ ), .B1(\keyboard/_0544_ ), .B2(\keyboard/_0431_ ), .ZN(\keyboard/_0545_ ) );
AOI21_X1 \keyboard/_0895_ ( .A(\keyboard/_0545_ ), .B1(\keyboard/_0431_ ), .B2(\keyboard/_0544_ ), .ZN(\keyboard/_0250_ ) );
AND2_X1 \keyboard/_0896_ ( .A1(\keyboard/_0524_ ), .A2(\keyboard/_0543_ ), .ZN(\keyboard/_0546_ ) );
AOI211_X2 \keyboard/_0897_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0546_ ), .C1(\keyboard/_0264_ ), .C2(\keyboard/_0544_ ), .ZN(\keyboard/_0251_ ) );
NOR2_X1 \keyboard/_0898_ ( .A1(\keyboard/_0522_ ), .A2(\keyboard/_0544_ ), .ZN(\keyboard/_0547_ ) );
AOI211_X2 \keyboard/_0899_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0547_ ), .C1(\keyboard/_0259_ ), .C2(\keyboard/_0544_ ), .ZN(\keyboard/_0252_ ) );
XNOR2_X2 \keyboard/_0900_ ( .A(\keyboard/_0512_ ), .B(\keyboard/_0526_ ), .ZN(\keyboard/_0548_ ) );
NOR2_X2 \keyboard/_0901_ ( .A1(\keyboard/_0548_ ), .A2(\keyboard/_0536_ ), .ZN(\keyboard/_0549_ ) );
AOI211_X2 \keyboard/_0902_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0549_ ), .C1(\keyboard/_0265_ ), .C2(\keyboard/_0536_ ), .ZN(\keyboard/_0254_ ) );
AND2_X4 \keyboard/_0903_ ( .A1(\keyboard/_0526_ ), .A2(\keyboard/_0755_ ), .ZN(\keyboard/_0550_ ) );
NOR2_X4 \keyboard/_0904_ ( .A1(\keyboard/_0526_ ), .A2(\keyboard/_0755_ ), .ZN(\keyboard/_0551_ ) );
NOR3_X4 \keyboard/_0905_ ( .A1(\keyboard/_0520_ ), .A2(\keyboard/_0550_ ), .A3(\keyboard/_0551_ ), .ZN(\keyboard/_0552_ ) );
AOI211_X2 \keyboard/_0906_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0552_ ), .C1(\keyboard/_0260_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0255_ ) );
AND2_X4 \keyboard/_0907_ ( .A1(\keyboard/_0754_ ), .A2(\keyboard/_0755_ ), .ZN(\keyboard/_0553_ ) );
OR2_X1 \keyboard/_0908_ ( .A1(\keyboard/_0553_ ), .A2(\keyboard/_0756_ ), .ZN(\keyboard/_0554_ ) );
NAND2_X1 \keyboard/_0909_ ( .A1(\keyboard/_0553_ ), .A2(\keyboard/_0756_ ), .ZN(\keyboard/_0555_ ) );
AOI21_X2 \keyboard/_0910_ ( .A(\keyboard/_0519_ ), .B1(\keyboard/_0554_ ), .B2(\keyboard/_0555_ ), .ZN(\keyboard/_0556_ ) );
AOI211_X2 \keyboard/_0911_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0556_ ), .C1(\keyboard/_0261_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0256_ ) );
CLKBUF_X1 \keyboard/_0912_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0557_ ) );
BUF_X2 \keyboard/_0913_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0558_ ) );
MUX2_X1 \keyboard/_0914_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0266_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0559_ ) );
AND4_X1 \keyboard/_0915_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0559_ ), .ZN(\keyboard/_0560_ ) );
AOI211_X2 \keyboard/_0916_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0560_ ), .C1(\keyboard/_0266_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0239_ ) );
MUX2_X1 \keyboard/_0917_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0268_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0561_ ) );
AND4_X1 \keyboard/_0918_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0561_ ), .ZN(\keyboard/_0562_ ) );
AOI211_X2 \keyboard/_0919_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0562_ ), .C1(\keyboard/_0268_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0240_ ) );
MUX2_X1 \keyboard/_0920_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0270_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0563_ ) );
AND4_X1 \keyboard/_0921_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0563_ ), .ZN(\keyboard/_0564_ ) );
AOI211_X2 \keyboard/_0922_ ( .A(\keyboard/_0501_ ), .B(\keyboard/_0564_ ), .C1(\keyboard/_0270_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0241_ ) );
CLKBUF_X1 \keyboard/_0923_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0565_ ) );
MUX2_X1 \keyboard/_0924_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0272_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0566_ ) );
AND4_X1 \keyboard/_0925_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0566_ ), .ZN(\keyboard/_0567_ ) );
AOI211_X2 \keyboard/_0926_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0567_ ), .C1(\keyboard/_0272_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0242_ ) );
MUX2_X1 \keyboard/_0927_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0274_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0568_ ) );
AND4_X1 \keyboard/_0928_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0568_ ), .ZN(\keyboard/_0569_ ) );
AOI211_X2 \keyboard/_0929_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0569_ ), .C1(\keyboard/_0274_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0243_ ) );
MUX2_X1 \keyboard/_0930_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0276_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0570_ ) );
AND4_X1 \keyboard/_0931_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0570_ ), .ZN(\keyboard/_0571_ ) );
AOI211_X2 \keyboard/_0932_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0571_ ), .C1(\keyboard/_0276_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0244_ ) );
MUX2_X1 \keyboard/_0933_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0278_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0572_ ) );
AND4_X1 \keyboard/_0934_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0572_ ), .ZN(\keyboard/_0573_ ) );
AOI211_X2 \keyboard/_0935_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0573_ ), .C1(\keyboard/_0278_ ), .C2(\keyboard/_0521_ ), .ZN(\keyboard/_0245_ ) );
MUX2_X1 \keyboard/_0936_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0280_ ), .S(\keyboard/_0555_ ), .Z(\keyboard/_0574_ ) );
AND4_X1 \keyboard/_0937_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0533_ ), .A4(\keyboard/_0574_ ), .ZN(\keyboard/_0575_ ) );
BUF_X32 \keyboard/_0938_ ( .A(\keyboard/_0520_ ), .Z(\keyboard/_0576_ ) );
AOI211_X2 \keyboard/_0939_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0575_ ), .C1(\keyboard/_0280_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0246_ ) );
CLKBUF_X1 \keyboard/_0940_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0577_ ) );
NAND2_X1 \keyboard/_0941_ ( .A1(\keyboard/_0550_ ), .A2(\keyboard/_0756_ ), .ZN(\keyboard/_0578_ ) );
MUX2_X1 \keyboard/_0942_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0282_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0579_ ) );
AND4_X1 \keyboard/_0943_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0579_ ), .ZN(\keyboard/_0580_ ) );
AOI211_X2 \keyboard/_0944_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0580_ ), .C1(\keyboard/_0282_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0231_ ) );
MUX2_X1 \keyboard/_0945_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0283_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0581_ ) );
AND4_X1 \keyboard/_0946_ ( .A1(\keyboard/_0557_ ), .A2(\keyboard/_0558_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0581_ ), .ZN(\keyboard/_0582_ ) );
AOI211_X2 \keyboard/_0947_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0582_ ), .C1(\keyboard/_0283_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0232_ ) );
CLKBUF_X1 \keyboard/_0948_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0583_ ) );
BUF_X2 \keyboard/_0949_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0584_ ) );
MUX2_X1 \keyboard/_0950_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0284_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0585_ ) );
AND4_X1 \keyboard/_0951_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0585_ ), .ZN(\keyboard/_0586_ ) );
AOI211_X2 \keyboard/_0952_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0586_ ), .C1(\keyboard/_0284_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0233_ ) );
MUX2_X1 \keyboard/_0953_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0285_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0587_ ) );
AND4_X1 \keyboard/_0954_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0587_ ), .ZN(\keyboard/_0588_ ) );
AOI211_X2 \keyboard/_0955_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0588_ ), .C1(\keyboard/_0285_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0234_ ) );
MUX2_X1 \keyboard/_0956_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0286_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0589_ ) );
AND4_X1 \keyboard/_0957_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0589_ ), .ZN(\keyboard/_0590_ ) );
AOI211_X2 \keyboard/_0958_ ( .A(\keyboard/_0565_ ), .B(\keyboard/_0590_ ), .C1(\keyboard/_0286_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0235_ ) );
CLKBUF_X1 \keyboard/_0959_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0591_ ) );
MUX2_X1 \keyboard/_0960_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0287_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0592_ ) );
AND4_X1 \keyboard/_0961_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0592_ ), .ZN(\keyboard/_0593_ ) );
AOI211_X2 \keyboard/_0962_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0593_ ), .C1(\keyboard/_0287_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0236_ ) );
MUX2_X1 \keyboard/_0963_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0288_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0594_ ) );
AND4_X1 \keyboard/_0964_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0594_ ), .ZN(\keyboard/_0595_ ) );
AOI211_X2 \keyboard/_0965_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0595_ ), .C1(\keyboard/_0288_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0237_ ) );
MUX2_X1 \keyboard/_0966_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0289_ ), .S(\keyboard/_0578_ ), .Z(\keyboard/_0596_ ) );
AND4_X1 \keyboard/_0967_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0596_ ), .ZN(\keyboard/_0597_ ) );
AOI211_X2 \keyboard/_0968_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0597_ ), .C1(\keyboard/_0289_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0238_ ) );
NAND2_X1 \keyboard/_0969_ ( .A1(\keyboard/_0551_ ), .A2(\keyboard/_0756_ ), .ZN(\keyboard/_0598_ ) );
MUX2_X1 \keyboard/_0970_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0290_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0599_ ) );
AND4_X1 \keyboard/_0971_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0599_ ), .ZN(\keyboard/_0600_ ) );
AOI211_X2 \keyboard/_0972_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0600_ ), .C1(\keyboard/_0290_ ), .C2(\keyboard/_0576_ ), .ZN(\keyboard/_0223_ ) );
MUX2_X1 \keyboard/_0973_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0291_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0601_ ) );
AND4_X1 \keyboard/_0974_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0577_ ), .A4(\keyboard/_0601_ ), .ZN(\keyboard/_0602_ ) );
BUF_X32 \keyboard/_0975_ ( .A(\keyboard/_0520_ ), .Z(\keyboard/_0603_ ) );
AOI211_X2 \keyboard/_0976_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0602_ ), .C1(\keyboard/_0291_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0224_ ) );
CLKBUF_X1 \keyboard/_0977_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0604_ ) );
MUX2_X1 \keyboard/_0978_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0292_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0605_ ) );
AND4_X1 \keyboard/_0979_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0605_ ), .ZN(\keyboard/_0606_ ) );
AOI211_X2 \keyboard/_0980_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0606_ ), .C1(\keyboard/_0292_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0225_ ) );
MUX2_X1 \keyboard/_0981_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0293_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0607_ ) );
AND4_X1 \keyboard/_0982_ ( .A1(\keyboard/_0583_ ), .A2(\keyboard/_0584_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0607_ ), .ZN(\keyboard/_0608_ ) );
AOI211_X2 \keyboard/_0983_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0608_ ), .C1(\keyboard/_0293_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0226_ ) );
CLKBUF_X1 \keyboard/_0984_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0609_ ) );
BUF_X2 \keyboard/_0985_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0610_ ) );
MUX2_X1 \keyboard/_0986_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0294_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0611_ ) );
AND4_X1 \keyboard/_0987_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0611_ ), .ZN(\keyboard/_0612_ ) );
AOI211_X2 \keyboard/_0988_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0612_ ), .C1(\keyboard/_0294_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0227_ ) );
MUX2_X1 \keyboard/_0989_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0295_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0613_ ) );
AND4_X1 \keyboard/_0990_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0613_ ), .ZN(\keyboard/_0614_ ) );
AOI211_X2 \keyboard/_0991_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0614_ ), .C1(\keyboard/_0295_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0228_ ) );
MUX2_X1 \keyboard/_0992_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0296_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0615_ ) );
AND4_X1 \keyboard/_0993_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0615_ ), .ZN(\keyboard/_0616_ ) );
AOI211_X2 \keyboard/_0994_ ( .A(\keyboard/_0591_ ), .B(\keyboard/_0616_ ), .C1(\keyboard/_0296_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0229_ ) );
CLKBUF_X1 \keyboard/_0995_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0617_ ) );
MUX2_X1 \keyboard/_0996_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0297_ ), .S(\keyboard/_0598_ ), .Z(\keyboard/_0618_ ) );
AND4_X1 \keyboard/_0997_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0618_ ), .ZN(\keyboard/_0619_ ) );
AOI211_X2 \keyboard/_0998_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0619_ ), .C1(\keyboard/_0297_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0230_ ) );
NOR2_X4 \keyboard/_0999_ ( .A1(\keyboard/_0754_ ), .A2(\keyboard/_0755_ ), .ZN(\keyboard/_0620_ ) );
NAND2_X1 \keyboard/_1000_ ( .A1(\keyboard/_0620_ ), .A2(\keyboard/_0756_ ), .ZN(\keyboard/_0621_ ) );
MUX2_X1 \keyboard/_1001_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0298_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0622_ ) );
AND4_X1 \keyboard/_1002_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0622_ ), .ZN(\keyboard/_0623_ ) );
AOI211_X2 \keyboard/_1003_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0623_ ), .C1(\keyboard/_0298_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0215_ ) );
MUX2_X1 \keyboard/_1004_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0299_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0624_ ) );
AND4_X1 \keyboard/_1005_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0624_ ), .ZN(\keyboard/_0625_ ) );
AOI211_X2 \keyboard/_1006_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0625_ ), .C1(\keyboard/_0299_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0216_ ) );
MUX2_X1 \keyboard/_1007_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0300_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0626_ ) );
AND4_X1 \keyboard/_1008_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0626_ ), .ZN(\keyboard/_0627_ ) );
AOI211_X2 \keyboard/_1009_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0627_ ), .C1(\keyboard/_0300_ ), .C2(\keyboard/_0603_ ), .ZN(\keyboard/_0217_ ) );
MUX2_X1 \keyboard/_1010_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0301_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0628_ ) );
AND4_X1 \keyboard/_1011_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0604_ ), .A4(\keyboard/_0628_ ), .ZN(\keyboard/_0629_ ) );
BUF_X32 \keyboard/_1012_ ( .A(\keyboard/_0520_ ), .Z(\keyboard/_0630_ ) );
AOI211_X2 \keyboard/_1013_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0629_ ), .C1(\keyboard/_0301_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0218_ ) );
CLKBUF_X1 \keyboard/_1014_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0631_ ) );
MUX2_X1 \keyboard/_1015_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0302_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0632_ ) );
AND4_X1 \keyboard/_1016_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0632_ ), .ZN(\keyboard/_0633_ ) );
AOI211_X2 \keyboard/_1017_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0633_ ), .C1(\keyboard/_0302_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0219_ ) );
MUX2_X1 \keyboard/_1018_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0303_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0634_ ) );
AND4_X1 \keyboard/_1019_ ( .A1(\keyboard/_0609_ ), .A2(\keyboard/_0610_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0634_ ), .ZN(\keyboard/_0635_ ) );
AOI211_X2 \keyboard/_1020_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0635_ ), .C1(\keyboard/_0303_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0220_ ) );
CLKBUF_X1 \keyboard/_1021_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0636_ ) );
BUF_X4 \keyboard/_1022_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0637_ ) );
MUX2_X1 \keyboard/_1023_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0304_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0638_ ) );
AND4_X1 \keyboard/_1024_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0638_ ), .ZN(\keyboard/_0639_ ) );
AOI211_X2 \keyboard/_1025_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0639_ ), .C1(\keyboard/_0304_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0221_ ) );
MUX2_X1 \keyboard/_1026_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0305_ ), .S(\keyboard/_0621_ ), .Z(\keyboard/_0640_ ) );
AND4_X1 \keyboard/_1027_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0640_ ), .ZN(\keyboard/_0641_ ) );
AOI211_X2 \keyboard/_1028_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0641_ ), .C1(\keyboard/_0305_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0222_ ) );
NAND2_X1 \keyboard/_1029_ ( .A1(\keyboard/_0553_ ), .A2(\keyboard/_0261_ ), .ZN(\keyboard/_0642_ ) );
MUX2_X1 \keyboard/_1030_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0306_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0643_ ) );
AND4_X1 \keyboard/_1031_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0643_ ), .ZN(\keyboard/_0644_ ) );
AOI211_X2 \keyboard/_1032_ ( .A(\keyboard/_0617_ ), .B(\keyboard/_0644_ ), .C1(\keyboard/_0306_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0207_ ) );
CLKBUF_X1 \keyboard/_1033_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0645_ ) );
MUX2_X1 \keyboard/_1034_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0307_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0646_ ) );
AND4_X1 \keyboard/_1035_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0646_ ), .ZN(\keyboard/_0647_ ) );
AOI211_X2 \keyboard/_1036_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0647_ ), .C1(\keyboard/_0307_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0208_ ) );
MUX2_X1 \keyboard/_1037_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0308_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0648_ ) );
AND4_X1 \keyboard/_1038_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0648_ ), .ZN(\keyboard/_0649_ ) );
AOI211_X2 \keyboard/_1039_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0649_ ), .C1(\keyboard/_0308_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0209_ ) );
MUX2_X1 \keyboard/_1040_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0309_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0650_ ) );
AND4_X1 \keyboard/_1041_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0650_ ), .ZN(\keyboard/_0651_ ) );
AOI211_X2 \keyboard/_1042_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0651_ ), .C1(\keyboard/_0309_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0210_ ) );
MUX2_X1 \keyboard/_1043_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0310_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0652_ ) );
AND4_X1 \keyboard/_1044_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0652_ ), .ZN(\keyboard/_0653_ ) );
AOI211_X2 \keyboard/_1045_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0653_ ), .C1(\keyboard/_0310_ ), .C2(\keyboard/_0630_ ), .ZN(\keyboard/_0211_ ) );
MUX2_X1 \keyboard/_1046_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0311_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0654_ ) );
AND4_X2 \keyboard/_1047_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0631_ ), .A4(\keyboard/_0654_ ), .ZN(\keyboard/_0655_ ) );
BUF_X8 \keyboard/_1048_ ( .A(\keyboard/_0519_ ), .Z(\keyboard/_0656_ ) );
AOI211_X2 \keyboard/_1049_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0655_ ), .C1(\keyboard/_0311_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0212_ ) );
CLKBUF_X1 \keyboard/_1050_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0657_ ) );
MUX2_X1 \keyboard/_1051_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0312_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0658_ ) );
AND4_X2 \keyboard/_1052_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0658_ ), .ZN(\keyboard/_0659_ ) );
AOI211_X2 \keyboard/_1053_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0659_ ), .C1(\keyboard/_0312_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0213_ ) );
MUX2_X1 \keyboard/_1054_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0313_ ), .S(\keyboard/_0642_ ), .Z(\keyboard/_0660_ ) );
AND4_X2 \keyboard/_1055_ ( .A1(\keyboard/_0636_ ), .A2(\keyboard/_0637_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0660_ ), .ZN(\keyboard/_0661_ ) );
AOI211_X2 \keyboard/_1056_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0661_ ), .C1(\keyboard/_0313_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0214_ ) );
CLKBUF_X1 \keyboard/_1057_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0662_ ) );
BUF_X4 \keyboard/_1058_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0663_ ) );
NAND2_X1 \keyboard/_1059_ ( .A1(\keyboard/_0550_ ), .A2(\keyboard/_0261_ ), .ZN(\keyboard/_0664_ ) );
MUX2_X1 \keyboard/_1060_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0314_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0665_ ) );
AND4_X2 \keyboard/_1061_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0665_ ), .ZN(\keyboard/_0666_ ) );
AOI211_X2 \keyboard/_1062_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0666_ ), .C1(\keyboard/_0314_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0199_ ) );
MUX2_X1 \keyboard/_1063_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0315_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0667_ ) );
AND4_X2 \keyboard/_1064_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0667_ ), .ZN(\keyboard/_0668_ ) );
AOI211_X2 \keyboard/_1065_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0668_ ), .C1(\keyboard/_0315_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0200_ ) );
MUX2_X1 \keyboard/_1066_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0316_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0669_ ) );
AND4_X2 \keyboard/_1067_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0669_ ), .ZN(\keyboard/_0670_ ) );
AOI211_X2 \keyboard/_1068_ ( .A(\keyboard/_0645_ ), .B(\keyboard/_0670_ ), .C1(\keyboard/_0316_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0201_ ) );
CLKBUF_X1 \keyboard/_1069_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0671_ ) );
MUX2_X1 \keyboard/_1070_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0317_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0672_ ) );
AND4_X2 \keyboard/_1071_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0672_ ), .ZN(\keyboard/_0673_ ) );
AOI211_X2 \keyboard/_1072_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0673_ ), .C1(\keyboard/_0317_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0202_ ) );
MUX2_X1 \keyboard/_1073_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0318_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0674_ ) );
AND4_X2 \keyboard/_1074_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0674_ ), .ZN(\keyboard/_0675_ ) );
AOI211_X2 \keyboard/_1075_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0675_ ), .C1(\keyboard/_0318_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0203_ ) );
MUX2_X1 \keyboard/_1076_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0319_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0676_ ) );
AND4_X2 \keyboard/_1077_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0676_ ), .ZN(\keyboard/_0677_ ) );
AOI211_X2 \keyboard/_1078_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0677_ ), .C1(\keyboard/_0319_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0204_ ) );
MUX2_X1 \keyboard/_1079_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0320_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0678_ ) );
AND4_X2 \keyboard/_1080_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0678_ ), .ZN(\keyboard/_0679_ ) );
AOI211_X2 \keyboard/_1081_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0679_ ), .C1(\keyboard/_0320_ ), .C2(\keyboard/_0656_ ), .ZN(\keyboard/_0205_ ) );
MUX2_X1 \keyboard/_1082_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0321_ ), .S(\keyboard/_0664_ ), .Z(\keyboard/_0680_ ) );
AND4_X2 \keyboard/_1083_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0657_ ), .A4(\keyboard/_0680_ ), .ZN(\keyboard/_0681_ ) );
BUF_X8 \keyboard/_1084_ ( .A(\keyboard/_0519_ ), .Z(\keyboard/_0682_ ) );
AOI211_X2 \keyboard/_1085_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0681_ ), .C1(\keyboard/_0321_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0206_ ) );
CLKBUF_X1 \keyboard/_1086_ ( .A(\keyboard/_0532_ ), .Z(\keyboard/_0683_ ) );
NAND2_X1 \keyboard/_1087_ ( .A1(\keyboard/_0551_ ), .A2(\keyboard/_0261_ ), .ZN(\keyboard/_0684_ ) );
MUX2_X1 \keyboard/_1088_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0322_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0685_ ) );
AND4_X2 \keyboard/_1089_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0685_ ), .ZN(\keyboard/_0686_ ) );
AOI211_X2 \keyboard/_1090_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0686_ ), .C1(\keyboard/_0322_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0191_ ) );
MUX2_X1 \keyboard/_1091_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0323_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0687_ ) );
AND4_X2 \keyboard/_1092_ ( .A1(\keyboard/_0662_ ), .A2(\keyboard/_0663_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0687_ ), .ZN(\keyboard/_0688_ ) );
AOI211_X2 \keyboard/_1093_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0688_ ), .C1(\keyboard/_0323_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0192_ ) );
CLKBUF_X1 \keyboard/_1094_ ( .A(\keyboard/_0511_ ), .Z(\keyboard/_0689_ ) );
BUF_X4 \keyboard/_1095_ ( .A(\keyboard/_0509_ ), .Z(\keyboard/_0690_ ) );
MUX2_X1 \keyboard/_1096_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0324_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0691_ ) );
AND4_X2 \keyboard/_1097_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0691_ ), .ZN(\keyboard/_0692_ ) );
AOI211_X2 \keyboard/_1098_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0692_ ), .C1(\keyboard/_0324_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0193_ ) );
MUX2_X1 \keyboard/_1099_ ( .A(\keyboard/_0273_ ), .B(\keyboard/_0325_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0693_ ) );
AND4_X2 \keyboard/_1100_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0693_ ), .ZN(\keyboard/_0694_ ) );
AOI211_X2 \keyboard/_1101_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0694_ ), .C1(\keyboard/_0325_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0194_ ) );
MUX2_X1 \keyboard/_1102_ ( .A(\keyboard/_0275_ ), .B(\keyboard/_0326_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0695_ ) );
AND4_X2 \keyboard/_1103_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0695_ ), .ZN(\keyboard/_0696_ ) );
AOI211_X2 \keyboard/_1104_ ( .A(\keyboard/_0671_ ), .B(\keyboard/_0696_ ), .C1(\keyboard/_0326_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0195_ ) );
CLKBUF_X1 \keyboard/_1105_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0697_ ) );
MUX2_X1 \keyboard/_1106_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0327_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0698_ ) );
AND4_X2 \keyboard/_1107_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0698_ ), .ZN(\keyboard/_0699_ ) );
AOI211_X2 \keyboard/_1108_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0699_ ), .C1(\keyboard/_0327_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0196_ ) );
MUX2_X1 \keyboard/_1109_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0328_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0700_ ) );
AND4_X2 \keyboard/_1110_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0700_ ), .ZN(\keyboard/_0701_ ) );
AOI211_X2 \keyboard/_1111_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0701_ ), .C1(\keyboard/_0328_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0197_ ) );
MUX2_X1 \keyboard/_1112_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0329_ ), .S(\keyboard/_0684_ ), .Z(\keyboard/_0702_ ) );
AND4_X2 \keyboard/_1113_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0702_ ), .ZN(\keyboard/_0703_ ) );
AOI211_X2 \keyboard/_1114_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0703_ ), .C1(\keyboard/_0329_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0198_ ) );
NAND2_X1 \keyboard/_1115_ ( .A1(\keyboard/_0620_ ), .A2(\keyboard/_0261_ ), .ZN(\keyboard/_0704_ ) );
MUX2_X1 \keyboard/_1116_ ( .A(\keyboard/_0267_ ), .B(\keyboard/_0330_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0705_ ) );
AND4_X2 \keyboard/_1117_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0705_ ), .ZN(\keyboard/_0706_ ) );
AOI211_X2 \keyboard/_1118_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0706_ ), .C1(\keyboard/_0330_ ), .C2(\keyboard/_0682_ ), .ZN(\keyboard/_0183_ ) );
MUX2_X1 \keyboard/_1119_ ( .A(\keyboard/_0269_ ), .B(\keyboard/_0331_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0707_ ) );
AND4_X2 \keyboard/_1120_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0683_ ), .A4(\keyboard/_0707_ ), .ZN(\keyboard/_0708_ ) );
AOI211_X2 \keyboard/_1121_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0708_ ), .C1(\keyboard/_0331_ ), .C2(\keyboard/_0520_ ), .ZN(\keyboard/_0184_ ) );
MUX2_X1 \keyboard/_1122_ ( .A(\keyboard/_0271_ ), .B(\keyboard/_0332_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0709_ ) );
AND4_X2 \keyboard/_1123_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0532_ ), .A4(\keyboard/_0709_ ), .ZN(\keyboard/_0710_ ) );
AOI211_X2 \keyboard/_1124_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0710_ ), .C1(\keyboard/_0332_ ), .C2(\keyboard/_0520_ ), .ZN(\keyboard/_0185_ ) );
NAND3_X4 \keyboard/_1125_ ( .A1(\keyboard/_0512_ ), .A2(\keyboard/_0517_ ), .A3(\keyboard/_0514_ ), .ZN(\keyboard/_0711_ ) );
NOR2_X2 \keyboard/_1126_ ( .A1(\keyboard/_0711_ ), .A2(\keyboard/_0704_ ), .ZN(\keyboard/_0712_ ) );
OAI21_X1 \keyboard/_1127_ ( .A(\keyboard/_0530_ ), .B1(\keyboard/_0712_ ), .B2(\keyboard/_0333_ ), .ZN(\keyboard/_0713_ ) );
NOR3_X1 \keyboard/_1128_ ( .A1(\keyboard/_0711_ ), .A2(\keyboard/_0273_ ), .A3(\keyboard/_0704_ ), .ZN(\keyboard/_0714_ ) );
NOR2_X1 \keyboard/_1129_ ( .A1(\keyboard/_0713_ ), .A2(\keyboard/_0714_ ), .ZN(\keyboard/_0715_ ) );
AOI211_X2 \keyboard/_1130_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0715_ ), .C1(\keyboard/_0333_ ), .C2(\keyboard/_0535_ ), .ZN(\keyboard/_0186_ ) );
OAI21_X1 \keyboard/_1131_ ( .A(\keyboard/_0530_ ), .B1(\keyboard/_0712_ ), .B2(\keyboard/_0334_ ), .ZN(\keyboard/_0716_ ) );
NOR3_X1 \keyboard/_1132_ ( .A1(\keyboard/_0711_ ), .A2(\keyboard/_0275_ ), .A3(\keyboard/_0704_ ), .ZN(\keyboard/_0717_ ) );
NOR2_X1 \keyboard/_1133_ ( .A1(\keyboard/_0716_ ), .A2(\keyboard/_0717_ ), .ZN(\keyboard/_0718_ ) );
AOI211_X2 \keyboard/_1134_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0718_ ), .C1(\keyboard/_0334_ ), .C2(\keyboard/_0535_ ), .ZN(\keyboard/_0187_ ) );
MUX2_X1 \keyboard/_1135_ ( .A(\keyboard/_0277_ ), .B(\keyboard/_0335_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0719_ ) );
AND4_X2 \keyboard/_1136_ ( .A1(\keyboard/_0689_ ), .A2(\keyboard/_0690_ ), .A3(\keyboard/_0532_ ), .A4(\keyboard/_0719_ ), .ZN(\keyboard/_0720_ ) );
AOI211_X2 \keyboard/_1137_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0720_ ), .C1(\keyboard/_0335_ ), .C2(\keyboard/_0520_ ), .ZN(\keyboard/_0188_ ) );
MUX2_X1 \keyboard/_1138_ ( .A(\keyboard/_0279_ ), .B(\keyboard/_0336_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0721_ ) );
AND4_X1 \keyboard/_1139_ ( .A1(\keyboard/_0511_ ), .A2(\keyboard/_0509_ ), .A3(\keyboard/_0532_ ), .A4(\keyboard/_0721_ ), .ZN(\keyboard/_0722_ ) );
AOI211_X2 \keyboard/_1140_ ( .A(\keyboard/_0697_ ), .B(\keyboard/_0722_ ), .C1(\keyboard/_0336_ ), .C2(\keyboard/_0520_ ), .ZN(\keyboard/_0189_ ) );
BUF_X8 \keyboard/_1141_ ( .A(\keyboard/_0500_ ), .Z(\keyboard/_0723_ ) );
MUX2_X1 \keyboard/_1142_ ( .A(\keyboard/_0281_ ), .B(\keyboard/_0337_ ), .S(\keyboard/_0704_ ), .Z(\keyboard/_0724_ ) );
AND4_X1 \keyboard/_1143_ ( .A1(\keyboard/_0511_ ), .A2(\keyboard/_0509_ ), .A3(\keyboard/_0532_ ), .A4(\keyboard/_0724_ ), .ZN(\keyboard/_0725_ ) );
AOI211_X2 \keyboard/_1144_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0725_ ), .C1(\keyboard/_0337_ ), .C2(\keyboard/_0520_ ), .ZN(\keyboard/_0190_ ) );
NOR3_X4 \keyboard/_1145_ ( .A1(\keyboard/_0535_ ), .A2(\keyboard/_0350_ ), .A3(\keyboard/_0351_ ), .ZN(\keyboard/_0726_ ) );
NOR2_X4 \keyboard/_1146_ ( .A1(\keyboard/_0352_ ), .A2(\keyboard/_0353_ ), .ZN(\keyboard/_0727_ ) );
AND3_X2 \keyboard/_1147_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0510_ ), .A3(\keyboard/_0727_ ), .ZN(\keyboard/_0728_ ) );
NAND2_X1 \keyboard/_1148_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0727_ ), .ZN(\keyboard/_0729_ ) );
AOI211_X2 \keyboard/_1149_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0728_ ), .C1(\keyboard/_0338_ ), .C2(\keyboard/_0729_ ), .ZN(\keyboard/_0169_ ) );
NAND3_X1 \keyboard/_1150_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0513_ ), .A3(\keyboard/_0727_ ), .ZN(\keyboard/_0730_ ) );
NOR2_X2 \keyboard/_1151_ ( .A1(\keyboard/_0730_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0731_ ) );
AOI211_X2 \keyboard/_1152_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0731_ ), .C1(\keyboard/_0267_ ), .C2(\keyboard/_0730_ ), .ZN(\keyboard/_0170_ ) );
NAND3_X1 \keyboard/_1153_ ( .A1(\keyboard/_0530_ ), .A2(\keyboard/_0514_ ), .A3(\keyboard/_0727_ ), .ZN(\keyboard/_0732_ ) );
NOR2_X1 \keyboard/_1154_ ( .A1(\keyboard/_0732_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0733_ ) );
AOI211_X2 \keyboard/_1155_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0733_ ), .C1(\keyboard/_0269_ ), .C2(\keyboard/_0732_ ), .ZN(\keyboard/_0171_ ) );
NAND3_X1 \keyboard/_1156_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0351_ ), .A3(\keyboard/_0727_ ), .ZN(\keyboard/_0734_ ) );
NOR2_X2 \keyboard/_1157_ ( .A1(\keyboard/_0734_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0735_ ) );
AOI211_X2 \keyboard/_1158_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0735_ ), .C1(\keyboard/_0271_ ), .C2(\keyboard/_0734_ ), .ZN(\keyboard/_0172_ ) );
AND2_X1 \keyboard/_1159_ ( .A1(\keyboard/_0516_ ), .A2(\keyboard/_0352_ ), .ZN(\keyboard/_0736_ ) );
AND3_X2 \keyboard/_1160_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0510_ ), .A3(\keyboard/_0736_ ), .ZN(\keyboard/_0737_ ) );
NAND2_X1 \keyboard/_1161_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0736_ ), .ZN(\keyboard/_0738_ ) );
AOI211_X2 \keyboard/_1162_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0737_ ), .C1(\keyboard/_0273_ ), .C2(\keyboard/_0738_ ), .ZN(\keyboard/_0173_ ) );
NAND3_X1 \keyboard/_1163_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0513_ ), .A3(\keyboard/_0736_ ), .ZN(\keyboard/_0739_ ) );
NOR2_X2 \keyboard/_1164_ ( .A1(\keyboard/_0739_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0740_ ) );
AOI211_X2 \keyboard/_1165_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0740_ ), .C1(\keyboard/_0275_ ), .C2(\keyboard/_0739_ ), .ZN(\keyboard/_0174_ ) );
NAND3_X1 \keyboard/_1166_ ( .A1(\keyboard/_0530_ ), .A2(\keyboard/_0736_ ), .A3(\keyboard/_0514_ ), .ZN(\keyboard/_0741_ ) );
NOR2_X1 \keyboard/_1167_ ( .A1(\keyboard/_0741_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0742_ ) );
AOI211_X2 \keyboard/_1168_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0742_ ), .C1(\keyboard/_0277_ ), .C2(\keyboard/_0741_ ), .ZN(\keyboard/_0175_ ) );
NAND3_X1 \keyboard/_1169_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0351_ ), .A3(\keyboard/_0736_ ), .ZN(\keyboard/_0743_ ) );
NOR2_X2 \keyboard/_1170_ ( .A1(\keyboard/_0743_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0744_ ) );
AOI211_X2 \keyboard/_1171_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0744_ ), .C1(\keyboard/_0279_ ), .C2(\keyboard/_0743_ ), .ZN(\keyboard/_0176_ ) );
AND3_X2 \keyboard/_1172_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0510_ ), .A3(\keyboard/_0517_ ), .ZN(\keyboard/_0745_ ) );
NAND2_X1 \keyboard/_1173_ ( .A1(\keyboard/_0726_ ), .A2(\keyboard/_0517_ ), .ZN(\keyboard/_0746_ ) );
AOI211_X2 \keyboard/_1174_ ( .A(\keyboard/_0723_ ), .B(\keyboard/_0745_ ), .C1(\keyboard/_0281_ ), .C2(\keyboard/_0746_ ), .ZN(\keyboard/_0177_ ) );
NAND3_X1 \keyboard/_1175_ ( .A1(\keyboard/_0531_ ), .A2(\keyboard/_0513_ ), .A3(\keyboard/_0517_ ), .ZN(\keyboard/_0747_ ) );
NOR2_X2 \keyboard/_1176_ ( .A1(\keyboard/_0747_ ), .A2(\keyboard/_0429_ ), .ZN(\keyboard/_0748_ ) );
AOI211_X2 \keyboard/_1177_ ( .A(\keyboard/_0500_ ), .B(\keyboard/_0748_ ), .C1(\keyboard/_0339_ ), .C2(\keyboard/_0747_ ), .ZN(\keyboard/_0178_ ) );
BUF_X1 \keyboard/_1178_ ( .A(io_ps2_clk ), .Z(\keyboard/_ps2_clk_sync_T_1[0] ) );
BUF_X1 \keyboard/_1179_ ( .A(\keyboard/_ps2_clk_sync_T_1[1] ), .Z(\keyboard/ps2_clk_sync[0] ) );
BUF_X1 \keyboard/_1180_ ( .A(\keyboard/_ps2_clk_sync_T_1[2] ), .Z(\keyboard/ps2_clk_sync[1] ) );
BUF_X1 \keyboard/_1181_ ( .A(\keyboard/r_ptr[1] ), .Z(\keyboard/_0751_ ) );
BUF_X1 \keyboard/_1182_ ( .A(\keyboard/r_ptr[0] ), .Z(\keyboard/_0750_ ) );
BUF_X1 \keyboard/_1183_ ( .A(\keyboard/r_ptr[2] ), .Z(\keyboard/_0752_ ) );
BUF_X1 \keyboard/_1184_ ( .A(\keyboard/_0088_ ), .Z(\keyboard/_0259_ ) );
BUF_X1 \keyboard/_1185_ ( .A(\keyboard/fifo_0[0] ), .Z(\keyboard/_0354_ ) );
BUF_X1 \keyboard/_1186_ ( .A(\keyboard/fifo_1[0] ), .Z(\keyboard/_0362_ ) );
BUF_X1 \keyboard/_1187_ ( .A(\keyboard/fifo_2[0] ), .Z(\keyboard/_0370_ ) );
BUF_X1 \keyboard/_1188_ ( .A(\keyboard/fifo_3[0] ), .Z(\keyboard/_0378_ ) );
BUF_X1 \keyboard/_1189_ ( .A(\keyboard/fifo_4[0] ), .Z(\keyboard/_0386_ ) );
BUF_X1 \keyboard/_1190_ ( .A(\keyboard/fifo_5[0] ), .Z(\keyboard/_0394_ ) );
BUF_X1 \keyboard/_1191_ ( .A(\keyboard/fifo_6[0] ), .Z(\keyboard/_0402_ ) );
BUF_X1 \keyboard/_1192_ ( .A(\keyboard/fifo_7[0] ), .Z(\keyboard/_0410_ ) );
BUF_X1 \keyboard/_1193_ ( .A(\keyboard/_0419_ ), .Z(\keyboard_io_data[0] ) );
BUF_X1 \keyboard/_1194_ ( .A(\keyboard/fifo_0[1] ), .Z(\keyboard/_0355_ ) );
BUF_X1 \keyboard/_1195_ ( .A(\keyboard/fifo_1[1] ), .Z(\keyboard/_0363_ ) );
BUF_X1 \keyboard/_1196_ ( .A(\keyboard/fifo_2[1] ), .Z(\keyboard/_0371_ ) );
BUF_X1 \keyboard/_1197_ ( .A(\keyboard/fifo_3[1] ), .Z(\keyboard/_0379_ ) );
BUF_X1 \keyboard/_1198_ ( .A(\keyboard/fifo_4[1] ), .Z(\keyboard/_0387_ ) );
BUF_X1 \keyboard/_1199_ ( .A(\keyboard/fifo_5[1] ), .Z(\keyboard/_0395_ ) );
BUF_X1 \keyboard/_1200_ ( .A(\keyboard/fifo_6[1] ), .Z(\keyboard/_0403_ ) );
BUF_X1 \keyboard/_1201_ ( .A(\keyboard/fifo_7[1] ), .Z(\keyboard/_0411_ ) );
BUF_X1 \keyboard/_1202_ ( .A(\keyboard/_0420_ ), .Z(\keyboard_io_data[1] ) );
BUF_X1 \keyboard/_1203_ ( .A(\keyboard/fifo_0[2] ), .Z(\keyboard/_0356_ ) );
BUF_X1 \keyboard/_1204_ ( .A(\keyboard/fifo_1[2] ), .Z(\keyboard/_0364_ ) );
BUF_X1 \keyboard/_1205_ ( .A(\keyboard/fifo_2[2] ), .Z(\keyboard/_0372_ ) );
BUF_X1 \keyboard/_1206_ ( .A(\keyboard/fifo_3[2] ), .Z(\keyboard/_0380_ ) );
BUF_X1 \keyboard/_1207_ ( .A(\keyboard/fifo_4[2] ), .Z(\keyboard/_0388_ ) );
BUF_X1 \keyboard/_1208_ ( .A(\keyboard/fifo_5[2] ), .Z(\keyboard/_0396_ ) );
BUF_X1 \keyboard/_1209_ ( .A(\keyboard/fifo_6[2] ), .Z(\keyboard/_0404_ ) );
BUF_X1 \keyboard/_1210_ ( .A(\keyboard/fifo_7[2] ), .Z(\keyboard/_0412_ ) );
BUF_X1 \keyboard/_1211_ ( .A(\keyboard/_0421_ ), .Z(\keyboard_io_data[2] ) );
BUF_X1 \keyboard/_1212_ ( .A(\keyboard/fifo_0[3] ), .Z(\keyboard/_0357_ ) );
BUF_X1 \keyboard/_1213_ ( .A(\keyboard/fifo_1[3] ), .Z(\keyboard/_0365_ ) );
BUF_X1 \keyboard/_1214_ ( .A(\keyboard/fifo_2[3] ), .Z(\keyboard/_0373_ ) );
BUF_X1 \keyboard/_1215_ ( .A(\keyboard/fifo_3[3] ), .Z(\keyboard/_0381_ ) );
BUF_X1 \keyboard/_1216_ ( .A(\keyboard/fifo_4[3] ), .Z(\keyboard/_0389_ ) );
BUF_X1 \keyboard/_1217_ ( .A(\keyboard/fifo_5[3] ), .Z(\keyboard/_0397_ ) );
BUF_X1 \keyboard/_1218_ ( .A(\keyboard/fifo_6[3] ), .Z(\keyboard/_0405_ ) );
BUF_X1 \keyboard/_1219_ ( .A(\keyboard/fifo_7[3] ), .Z(\keyboard/_0413_ ) );
BUF_X1 \keyboard/_1220_ ( .A(\keyboard/_0422_ ), .Z(\keyboard_io_data[3] ) );
BUF_X1 \keyboard/_1221_ ( .A(\keyboard/fifo_0[4] ), .Z(\keyboard/_0358_ ) );
BUF_X1 \keyboard/_1222_ ( .A(\keyboard/fifo_1[4] ), .Z(\keyboard/_0366_ ) );
BUF_X1 \keyboard/_1223_ ( .A(\keyboard/fifo_2[4] ), .Z(\keyboard/_0374_ ) );
BUF_X1 \keyboard/_1224_ ( .A(\keyboard/fifo_3[4] ), .Z(\keyboard/_0382_ ) );
BUF_X1 \keyboard/_1225_ ( .A(\keyboard/fifo_4[4] ), .Z(\keyboard/_0390_ ) );
BUF_X1 \keyboard/_1226_ ( .A(\keyboard/fifo_5[4] ), .Z(\keyboard/_0398_ ) );
BUF_X1 \keyboard/_1227_ ( .A(\keyboard/fifo_6[4] ), .Z(\keyboard/_0406_ ) );
BUF_X1 \keyboard/_1228_ ( .A(\keyboard/fifo_7[4] ), .Z(\keyboard/_0414_ ) );
BUF_X1 \keyboard/_1229_ ( .A(\keyboard/_0423_ ), .Z(\keyboard_io_data[4] ) );
BUF_X1 \keyboard/_1230_ ( .A(\keyboard/fifo_0[5] ), .Z(\keyboard/_0359_ ) );
BUF_X1 \keyboard/_1231_ ( .A(\keyboard/fifo_1[5] ), .Z(\keyboard/_0367_ ) );
BUF_X1 \keyboard/_1232_ ( .A(\keyboard/fifo_2[5] ), .Z(\keyboard/_0375_ ) );
BUF_X1 \keyboard/_1233_ ( .A(\keyboard/fifo_3[5] ), .Z(\keyboard/_0383_ ) );
BUF_X1 \keyboard/_1234_ ( .A(\keyboard/fifo_4[5] ), .Z(\keyboard/_0391_ ) );
BUF_X1 \keyboard/_1235_ ( .A(\keyboard/fifo_5[5] ), .Z(\keyboard/_0399_ ) );
BUF_X1 \keyboard/_1236_ ( .A(\keyboard/fifo_6[5] ), .Z(\keyboard/_0407_ ) );
BUF_X1 \keyboard/_1237_ ( .A(\keyboard/fifo_7[5] ), .Z(\keyboard/_0415_ ) );
BUF_X1 \keyboard/_1238_ ( .A(\keyboard/_0424_ ), .Z(\keyboard_io_data[5] ) );
BUF_X1 \keyboard/_1239_ ( .A(\keyboard/fifo_0[6] ), .Z(\keyboard/_0360_ ) );
BUF_X1 \keyboard/_1240_ ( .A(\keyboard/fifo_1[6] ), .Z(\keyboard/_0368_ ) );
BUF_X1 \keyboard/_1241_ ( .A(\keyboard/fifo_2[6] ), .Z(\keyboard/_0376_ ) );
BUF_X1 \keyboard/_1242_ ( .A(\keyboard/fifo_3[6] ), .Z(\keyboard/_0384_ ) );
BUF_X1 \keyboard/_1243_ ( .A(\keyboard/fifo_4[6] ), .Z(\keyboard/_0392_ ) );
BUF_X1 \keyboard/_1244_ ( .A(\keyboard/fifo_5[6] ), .Z(\keyboard/_0400_ ) );
BUF_X1 \keyboard/_1245_ ( .A(\keyboard/fifo_6[6] ), .Z(\keyboard/_0408_ ) );
BUF_X1 \keyboard/_1246_ ( .A(\keyboard/fifo_7[6] ), .Z(\keyboard/_0416_ ) );
BUF_X1 \keyboard/_1247_ ( .A(\keyboard/_0425_ ), .Z(\keyboard_io_data[6] ) );
BUF_X1 \keyboard/_1248_ ( .A(\keyboard/fifo_0[7] ), .Z(\keyboard/_0361_ ) );
BUF_X1 \keyboard/_1249_ ( .A(\keyboard/fifo_1[7] ), .Z(\keyboard/_0369_ ) );
BUF_X1 \keyboard/_1250_ ( .A(\keyboard/fifo_2[7] ), .Z(\keyboard/_0377_ ) );
BUF_X1 \keyboard/_1251_ ( .A(\keyboard/fifo_3[7] ), .Z(\keyboard/_0385_ ) );
BUF_X1 \keyboard/_1252_ ( .A(\keyboard/fifo_4[7] ), .Z(\keyboard/_0393_ ) );
BUF_X1 \keyboard/_1253_ ( .A(\keyboard/fifo_5[7] ), .Z(\keyboard/_0401_ ) );
BUF_X1 \keyboard/_1254_ ( .A(\keyboard/fifo_6[7] ), .Z(\keyboard/_0409_ ) );
BUF_X1 \keyboard/_1255_ ( .A(\keyboard/fifo_7[7] ), .Z(\keyboard/_0417_ ) );
BUF_X1 \keyboard/_1256_ ( .A(\keyboard/_0426_ ), .Z(\keyboard_io_data[7] ) );
BUF_X1 \keyboard/_1257_ ( .A(io_ps2_clk ), .Z(\keyboard/_0428_ ) );
BUF_X1 \keyboard/_1258_ ( .A(reset ), .Z(\keyboard/_0753_ ) );
BUF_X1 \keyboard/_1259_ ( .A(\keyboard/_0247_ ), .Z(\keyboard/_0078_ ) );
BUF_X1 \keyboard/_1260_ ( .A(\keyboard/_ps2_clk_sync_T_1[1] ), .Z(\keyboard/_0257_ ) );
BUF_X1 \keyboard/_1261_ ( .A(\keyboard/_0248_ ), .Z(\keyboard/_0079_ ) );
BUF_X1 \keyboard/_1262_ ( .A(\keyboard/_ps2_clk_sync_T_1[2] ), .Z(\keyboard/_0258_ ) );
BUF_X1 \keyboard/_1263_ ( .A(\keyboard/_0249_ ), .Z(\keyboard/_0080_ ) );
BUF_X1 \keyboard/_1264_ ( .A(keyboard_io_nextdata_n ), .Z(\keyboard/_0427_ ) );
BUF_X1 \keyboard/_1265_ ( .A(keyboard_io_ready ), .Z(\keyboard/_0430_ ) );
BUF_X1 \keyboard/_1266_ ( .A(\keyboard/w_ptr[0] ), .Z(\keyboard/_0754_ ) );
BUF_X1 \keyboard/_1267_ ( .A(\keyboard/_0089_ ), .Z(\keyboard/_0260_ ) );
BUF_X1 \keyboard/_1268_ ( .A(\keyboard/_0090_ ), .Z(\keyboard/_0261_ ) );
BUF_X1 \keyboard/_1269_ ( .A(\keyboard/ps2_clk_sync[2] ), .Z(\keyboard/_0749_ ) );
BUF_X1 \keyboard/_1270_ ( .A(io_ps2_data ), .Z(\keyboard/_0429_ ) );
BUF_X1 \keyboard/_1271_ ( .A(\keyboard/buffer[0] ), .Z(\keyboard/_0340_ ) );
BUF_X1 \keyboard/_1272_ ( .A(\keyboard/buffer[2] ), .Z(\keyboard/_0342_ ) );
BUF_X1 \keyboard/_1273_ ( .A(\keyboard/buffer[1] ), .Z(\keyboard/_0341_ ) );
BUF_X1 \keyboard/_1274_ ( .A(\keyboard/buffer[4] ), .Z(\keyboard/_0344_ ) );
BUF_X1 \keyboard/_1275_ ( .A(\keyboard/buffer[3] ), .Z(\keyboard/_0343_ ) );
BUF_X1 \keyboard/_1276_ ( .A(\keyboard/buffer[6] ), .Z(\keyboard/_0346_ ) );
BUF_X1 \keyboard/_1277_ ( .A(\keyboard/buffer[5] ), .Z(\keyboard/_0345_ ) );
BUF_X1 \keyboard/_1278_ ( .A(\keyboard/buffer[8] ), .Z(\keyboard/_0348_ ) );
BUF_X1 \keyboard/_1279_ ( .A(\keyboard/buffer[7] ), .Z(\keyboard/_0347_ ) );
BUF_X1 \keyboard/_1280_ ( .A(\keyboard/buffer[9] ), .Z(\keyboard/_0349_ ) );
BUF_X1 \keyboard/_1281_ ( .A(\keyboard/count[0] ), .Z(\keyboard/_0350_ ) );
BUF_X1 \keyboard/_1282_ ( .A(\keyboard/count[1] ), .Z(\keyboard/_0351_ ) );
BUF_X1 \keyboard/_1283_ ( .A(\keyboard/count[2] ), .Z(\keyboard/_0352_ ) );
BUF_X1 \keyboard/_1284_ ( .A(\keyboard/count[3] ), .Z(\keyboard/_0353_ ) );
BUF_X1 \keyboard/_1285_ ( .A(io_clrn ), .Z(\keyboard/_0418_ ) );
BUF_X1 \keyboard/_1286_ ( .A(\keyboard/_0253_ ), .Z(\keyboard/_0084_ ) );
BUF_X1 \keyboard/_1287_ ( .A(\keyboard/_0091_ ), .Z(\keyboard/_0262_ ) );
BUF_X1 \keyboard/_1288_ ( .A(\keyboard/_0179_ ), .Z(\keyboard/_0010_ ) );
BUF_X1 \keyboard/_1289_ ( .A(\keyboard/_0180_ ), .Z(\keyboard/_0011_ ) );
BUF_X1 \keyboard/_1290_ ( .A(\keyboard/_0181_ ), .Z(\keyboard/_0012_ ) );
BUF_X1 \keyboard/_1291_ ( .A(\keyboard/_0092_ ), .Z(\keyboard/_0263_ ) );
BUF_X1 \keyboard/_1292_ ( .A(\keyboard/_0182_ ), .Z(\keyboard/_0013_ ) );
BUF_X1 \keyboard/_1293_ ( .A(\keyboard/_0250_ ), .Z(\keyboard/_0081_ ) );
BUF_X1 \keyboard/_1294_ ( .A(\keyboard/_0093_ ), .Z(\keyboard/_0264_ ) );
BUF_X1 \keyboard/_1295_ ( .A(\keyboard/_0251_ ), .Z(\keyboard/_0082_ ) );
BUF_X1 \keyboard/_1296_ ( .A(\keyboard/_0252_ ), .Z(\keyboard/_0083_ ) );
BUF_X1 \keyboard/_1297_ ( .A(\keyboard/_0094_ ), .Z(\keyboard/_0265_ ) );
BUF_X1 \keyboard/_1298_ ( .A(\keyboard/_0254_ ), .Z(\keyboard/_0085_ ) );
BUF_X1 \keyboard/_1299_ ( .A(\keyboard/w_ptr[1] ), .Z(\keyboard/_0755_ ) );
BUF_X1 \keyboard/_1300_ ( .A(\keyboard/_0255_ ), .Z(\keyboard/_0086_ ) );
BUF_X1 \keyboard/_1301_ ( .A(\keyboard/w_ptr[2] ), .Z(\keyboard/_0756_ ) );
BUF_X1 \keyboard/_1302_ ( .A(\keyboard/_0256_ ), .Z(\keyboard/_0087_ ) );
BUF_X1 \keyboard/_1303_ ( .A(\keyboard/_0095_ ), .Z(\keyboard/_0266_ ) );
BUF_X1 \keyboard/_1304_ ( .A(\keyboard/_0096_ ), .Z(\keyboard/_0267_ ) );
BUF_X1 \keyboard/_1305_ ( .A(\keyboard/_0239_ ), .Z(\keyboard/_0070_ ) );
BUF_X1 \keyboard/_1306_ ( .A(\keyboard/_0097_ ), .Z(\keyboard/_0268_ ) );
BUF_X1 \keyboard/_1307_ ( .A(\keyboard/_0098_ ), .Z(\keyboard/_0269_ ) );
BUF_X1 \keyboard/_1308_ ( .A(\keyboard/_0240_ ), .Z(\keyboard/_0071_ ) );
BUF_X1 \keyboard/_1309_ ( .A(\keyboard/_0099_ ), .Z(\keyboard/_0270_ ) );
BUF_X1 \keyboard/_1310_ ( .A(\keyboard/_0100_ ), .Z(\keyboard/_0271_ ) );
BUF_X1 \keyboard/_1311_ ( .A(\keyboard/_0241_ ), .Z(\keyboard/_0072_ ) );
BUF_X1 \keyboard/_1312_ ( .A(\keyboard/_0101_ ), .Z(\keyboard/_0272_ ) );
BUF_X1 \keyboard/_1313_ ( .A(\keyboard/_0102_ ), .Z(\keyboard/_0273_ ) );
BUF_X1 \keyboard/_1314_ ( .A(\keyboard/_0242_ ), .Z(\keyboard/_0073_ ) );
BUF_X1 \keyboard/_1315_ ( .A(\keyboard/_0103_ ), .Z(\keyboard/_0274_ ) );
BUF_X1 \keyboard/_1316_ ( .A(\keyboard/_0104_ ), .Z(\keyboard/_0275_ ) );
BUF_X1 \keyboard/_1317_ ( .A(\keyboard/_0243_ ), .Z(\keyboard/_0074_ ) );
BUF_X1 \keyboard/_1318_ ( .A(\keyboard/_0105_ ), .Z(\keyboard/_0276_ ) );
BUF_X1 \keyboard/_1319_ ( .A(\keyboard/_0106_ ), .Z(\keyboard/_0277_ ) );
BUF_X1 \keyboard/_1320_ ( .A(\keyboard/_0244_ ), .Z(\keyboard/_0075_ ) );
BUF_X1 \keyboard/_1321_ ( .A(\keyboard/_0107_ ), .Z(\keyboard/_0278_ ) );
BUF_X1 \keyboard/_1322_ ( .A(\keyboard/_0108_ ), .Z(\keyboard/_0279_ ) );
BUF_X1 \keyboard/_1323_ ( .A(\keyboard/_0245_ ), .Z(\keyboard/_0076_ ) );
BUF_X1 \keyboard/_1324_ ( .A(\keyboard/_0109_ ), .Z(\keyboard/_0280_ ) );
BUF_X1 \keyboard/_1325_ ( .A(\keyboard/_0110_ ), .Z(\keyboard/_0281_ ) );
BUF_X1 \keyboard/_1326_ ( .A(\keyboard/_0246_ ), .Z(\keyboard/_0077_ ) );
BUF_X1 \keyboard/_1327_ ( .A(\keyboard/_0111_ ), .Z(\keyboard/_0282_ ) );
BUF_X1 \keyboard/_1328_ ( .A(\keyboard/_0231_ ), .Z(\keyboard/_0062_ ) );
BUF_X1 \keyboard/_1329_ ( .A(\keyboard/_0112_ ), .Z(\keyboard/_0283_ ) );
BUF_X1 \keyboard/_1330_ ( .A(\keyboard/_0232_ ), .Z(\keyboard/_0063_ ) );
BUF_X1 \keyboard/_1331_ ( .A(\keyboard/_0113_ ), .Z(\keyboard/_0284_ ) );
BUF_X1 \keyboard/_1332_ ( .A(\keyboard/_0233_ ), .Z(\keyboard/_0064_ ) );
BUF_X1 \keyboard/_1333_ ( .A(\keyboard/_0114_ ), .Z(\keyboard/_0285_ ) );
BUF_X1 \keyboard/_1334_ ( .A(\keyboard/_0234_ ), .Z(\keyboard/_0065_ ) );
BUF_X1 \keyboard/_1335_ ( .A(\keyboard/_0115_ ), .Z(\keyboard/_0286_ ) );
BUF_X1 \keyboard/_1336_ ( .A(\keyboard/_0235_ ), .Z(\keyboard/_0066_ ) );
BUF_X1 \keyboard/_1337_ ( .A(\keyboard/_0116_ ), .Z(\keyboard/_0287_ ) );
BUF_X1 \keyboard/_1338_ ( .A(\keyboard/_0236_ ), .Z(\keyboard/_0067_ ) );
BUF_X1 \keyboard/_1339_ ( .A(\keyboard/_0117_ ), .Z(\keyboard/_0288_ ) );
BUF_X1 \keyboard/_1340_ ( .A(\keyboard/_0237_ ), .Z(\keyboard/_0068_ ) );
BUF_X1 \keyboard/_1341_ ( .A(\keyboard/_0118_ ), .Z(\keyboard/_0289_ ) );
BUF_X1 \keyboard/_1342_ ( .A(\keyboard/_0238_ ), .Z(\keyboard/_0069_ ) );
BUF_X1 \keyboard/_1343_ ( .A(\keyboard/_0119_ ), .Z(\keyboard/_0290_ ) );
BUF_X1 \keyboard/_1344_ ( .A(\keyboard/_0223_ ), .Z(\keyboard/_0054_ ) );
BUF_X1 \keyboard/_1345_ ( .A(\keyboard/_0120_ ), .Z(\keyboard/_0291_ ) );
BUF_X1 \keyboard/_1346_ ( .A(\keyboard/_0224_ ), .Z(\keyboard/_0055_ ) );
BUF_X1 \keyboard/_1347_ ( .A(\keyboard/_0121_ ), .Z(\keyboard/_0292_ ) );
BUF_X1 \keyboard/_1348_ ( .A(\keyboard/_0225_ ), .Z(\keyboard/_0056_ ) );
BUF_X1 \keyboard/_1349_ ( .A(\keyboard/_0122_ ), .Z(\keyboard/_0293_ ) );
BUF_X1 \keyboard/_1350_ ( .A(\keyboard/_0226_ ), .Z(\keyboard/_0057_ ) );
BUF_X1 \keyboard/_1351_ ( .A(\keyboard/_0123_ ), .Z(\keyboard/_0294_ ) );
BUF_X1 \keyboard/_1352_ ( .A(\keyboard/_0227_ ), .Z(\keyboard/_0058_ ) );
BUF_X1 \keyboard/_1353_ ( .A(\keyboard/_0124_ ), .Z(\keyboard/_0295_ ) );
BUF_X1 \keyboard/_1354_ ( .A(\keyboard/_0228_ ), .Z(\keyboard/_0059_ ) );
BUF_X1 \keyboard/_1355_ ( .A(\keyboard/_0125_ ), .Z(\keyboard/_0296_ ) );
BUF_X1 \keyboard/_1356_ ( .A(\keyboard/_0229_ ), .Z(\keyboard/_0060_ ) );
BUF_X1 \keyboard/_1357_ ( .A(\keyboard/_0126_ ), .Z(\keyboard/_0297_ ) );
BUF_X1 \keyboard/_1358_ ( .A(\keyboard/_0230_ ), .Z(\keyboard/_0061_ ) );
BUF_X1 \keyboard/_1359_ ( .A(\keyboard/_0127_ ), .Z(\keyboard/_0298_ ) );
BUF_X1 \keyboard/_1360_ ( .A(\keyboard/_0215_ ), .Z(\keyboard/_0046_ ) );
BUF_X1 \keyboard/_1361_ ( .A(\keyboard/_0128_ ), .Z(\keyboard/_0299_ ) );
BUF_X1 \keyboard/_1362_ ( .A(\keyboard/_0216_ ), .Z(\keyboard/_0047_ ) );
BUF_X1 \keyboard/_1363_ ( .A(\keyboard/_0129_ ), .Z(\keyboard/_0300_ ) );
BUF_X1 \keyboard/_1364_ ( .A(\keyboard/_0217_ ), .Z(\keyboard/_0048_ ) );
BUF_X1 \keyboard/_1365_ ( .A(\keyboard/_0130_ ), .Z(\keyboard/_0301_ ) );
BUF_X1 \keyboard/_1366_ ( .A(\keyboard/_0218_ ), .Z(\keyboard/_0049_ ) );
BUF_X1 \keyboard/_1367_ ( .A(\keyboard/_0131_ ), .Z(\keyboard/_0302_ ) );
BUF_X1 \keyboard/_1368_ ( .A(\keyboard/_0219_ ), .Z(\keyboard/_0050_ ) );
BUF_X1 \keyboard/_1369_ ( .A(\keyboard/_0132_ ), .Z(\keyboard/_0303_ ) );
BUF_X1 \keyboard/_1370_ ( .A(\keyboard/_0220_ ), .Z(\keyboard/_0051_ ) );
BUF_X1 \keyboard/_1371_ ( .A(\keyboard/_0133_ ), .Z(\keyboard/_0304_ ) );
BUF_X1 \keyboard/_1372_ ( .A(\keyboard/_0221_ ), .Z(\keyboard/_0052_ ) );
BUF_X1 \keyboard/_1373_ ( .A(\keyboard/_0134_ ), .Z(\keyboard/_0305_ ) );
BUF_X1 \keyboard/_1374_ ( .A(\keyboard/_0222_ ), .Z(\keyboard/_0053_ ) );
BUF_X1 \keyboard/_1375_ ( .A(\keyboard/_0135_ ), .Z(\keyboard/_0306_ ) );
BUF_X1 \keyboard/_1376_ ( .A(\keyboard/_0207_ ), .Z(\keyboard/_0038_ ) );
BUF_X1 \keyboard/_1377_ ( .A(\keyboard/_0136_ ), .Z(\keyboard/_0307_ ) );
BUF_X1 \keyboard/_1378_ ( .A(\keyboard/_0208_ ), .Z(\keyboard/_0039_ ) );
BUF_X1 \keyboard/_1379_ ( .A(\keyboard/_0137_ ), .Z(\keyboard/_0308_ ) );
BUF_X1 \keyboard/_1380_ ( .A(\keyboard/_0209_ ), .Z(\keyboard/_0040_ ) );
BUF_X1 \keyboard/_1381_ ( .A(\keyboard/_0138_ ), .Z(\keyboard/_0309_ ) );
BUF_X1 \keyboard/_1382_ ( .A(\keyboard/_0210_ ), .Z(\keyboard/_0041_ ) );
BUF_X1 \keyboard/_1383_ ( .A(\keyboard/_0139_ ), .Z(\keyboard/_0310_ ) );
BUF_X1 \keyboard/_1384_ ( .A(\keyboard/_0211_ ), .Z(\keyboard/_0042_ ) );
BUF_X1 \keyboard/_1385_ ( .A(\keyboard/_0140_ ), .Z(\keyboard/_0311_ ) );
BUF_X1 \keyboard/_1386_ ( .A(\keyboard/_0212_ ), .Z(\keyboard/_0043_ ) );
BUF_X1 \keyboard/_1387_ ( .A(\keyboard/_0141_ ), .Z(\keyboard/_0312_ ) );
BUF_X1 \keyboard/_1388_ ( .A(\keyboard/_0213_ ), .Z(\keyboard/_0044_ ) );
BUF_X1 \keyboard/_1389_ ( .A(\keyboard/_0142_ ), .Z(\keyboard/_0313_ ) );
BUF_X1 \keyboard/_1390_ ( .A(\keyboard/_0214_ ), .Z(\keyboard/_0045_ ) );
BUF_X1 \keyboard/_1391_ ( .A(\keyboard/_0143_ ), .Z(\keyboard/_0314_ ) );
BUF_X1 \keyboard/_1392_ ( .A(\keyboard/_0199_ ), .Z(\keyboard/_0030_ ) );
BUF_X1 \keyboard/_1393_ ( .A(\keyboard/_0144_ ), .Z(\keyboard/_0315_ ) );
BUF_X1 \keyboard/_1394_ ( .A(\keyboard/_0200_ ), .Z(\keyboard/_0031_ ) );
BUF_X1 \keyboard/_1395_ ( .A(\keyboard/_0145_ ), .Z(\keyboard/_0316_ ) );
BUF_X1 \keyboard/_1396_ ( .A(\keyboard/_0201_ ), .Z(\keyboard/_0032_ ) );
BUF_X1 \keyboard/_1397_ ( .A(\keyboard/_0146_ ), .Z(\keyboard/_0317_ ) );
BUF_X1 \keyboard/_1398_ ( .A(\keyboard/_0202_ ), .Z(\keyboard/_0033_ ) );
BUF_X1 \keyboard/_1399_ ( .A(\keyboard/_0147_ ), .Z(\keyboard/_0318_ ) );
BUF_X1 \keyboard/_1400_ ( .A(\keyboard/_0203_ ), .Z(\keyboard/_0034_ ) );
BUF_X1 \keyboard/_1401_ ( .A(\keyboard/_0148_ ), .Z(\keyboard/_0319_ ) );
BUF_X1 \keyboard/_1402_ ( .A(\keyboard/_0204_ ), .Z(\keyboard/_0035_ ) );
BUF_X1 \keyboard/_1403_ ( .A(\keyboard/_0149_ ), .Z(\keyboard/_0320_ ) );
BUF_X1 \keyboard/_1404_ ( .A(\keyboard/_0205_ ), .Z(\keyboard/_0036_ ) );
BUF_X1 \keyboard/_1405_ ( .A(\keyboard/_0150_ ), .Z(\keyboard/_0321_ ) );
BUF_X1 \keyboard/_1406_ ( .A(\keyboard/_0206_ ), .Z(\keyboard/_0037_ ) );
BUF_X1 \keyboard/_1407_ ( .A(\keyboard/_0151_ ), .Z(\keyboard/_0322_ ) );
BUF_X1 \keyboard/_1408_ ( .A(\keyboard/_0191_ ), .Z(\keyboard/_0022_ ) );
BUF_X1 \keyboard/_1409_ ( .A(\keyboard/_0152_ ), .Z(\keyboard/_0323_ ) );
BUF_X1 \keyboard/_1410_ ( .A(\keyboard/_0192_ ), .Z(\keyboard/_0023_ ) );
BUF_X1 \keyboard/_1411_ ( .A(\keyboard/_0153_ ), .Z(\keyboard/_0324_ ) );
BUF_X1 \keyboard/_1412_ ( .A(\keyboard/_0193_ ), .Z(\keyboard/_0024_ ) );
BUF_X1 \keyboard/_1413_ ( .A(\keyboard/_0154_ ), .Z(\keyboard/_0325_ ) );
BUF_X1 \keyboard/_1414_ ( .A(\keyboard/_0194_ ), .Z(\keyboard/_0025_ ) );
BUF_X1 \keyboard/_1415_ ( .A(\keyboard/_0155_ ), .Z(\keyboard/_0326_ ) );
BUF_X1 \keyboard/_1416_ ( .A(\keyboard/_0195_ ), .Z(\keyboard/_0026_ ) );
BUF_X1 \keyboard/_1417_ ( .A(\keyboard/_0156_ ), .Z(\keyboard/_0327_ ) );
BUF_X1 \keyboard/_1418_ ( .A(\keyboard/_0196_ ), .Z(\keyboard/_0027_ ) );
BUF_X1 \keyboard/_1419_ ( .A(\keyboard/_0157_ ), .Z(\keyboard/_0328_ ) );
BUF_X1 \keyboard/_1420_ ( .A(\keyboard/_0197_ ), .Z(\keyboard/_0028_ ) );
BUF_X1 \keyboard/_1421_ ( .A(\keyboard/_0158_ ), .Z(\keyboard/_0329_ ) );
BUF_X1 \keyboard/_1422_ ( .A(\keyboard/_0198_ ), .Z(\keyboard/_0029_ ) );
BUF_X1 \keyboard/_1423_ ( .A(\keyboard/_0159_ ), .Z(\keyboard/_0330_ ) );
BUF_X1 \keyboard/_1424_ ( .A(\keyboard/_0183_ ), .Z(\keyboard/_0014_ ) );
BUF_X1 \keyboard/_1425_ ( .A(\keyboard/_0160_ ), .Z(\keyboard/_0331_ ) );
BUF_X1 \keyboard/_1426_ ( .A(\keyboard/_0184_ ), .Z(\keyboard/_0015_ ) );
BUF_X1 \keyboard/_1427_ ( .A(\keyboard/_0161_ ), .Z(\keyboard/_0332_ ) );
BUF_X1 \keyboard/_1428_ ( .A(\keyboard/_0185_ ), .Z(\keyboard/_0016_ ) );
BUF_X1 \keyboard/_1429_ ( .A(\keyboard/_0162_ ), .Z(\keyboard/_0333_ ) );
BUF_X1 \keyboard/_1430_ ( .A(\keyboard/_0186_ ), .Z(\keyboard/_0017_ ) );
BUF_X1 \keyboard/_1431_ ( .A(\keyboard/_0163_ ), .Z(\keyboard/_0334_ ) );
BUF_X1 \keyboard/_1432_ ( .A(\keyboard/_0187_ ), .Z(\keyboard/_0018_ ) );
BUF_X1 \keyboard/_1433_ ( .A(\keyboard/_0164_ ), .Z(\keyboard/_0335_ ) );
BUF_X1 \keyboard/_1434_ ( .A(\keyboard/_0188_ ), .Z(\keyboard/_0019_ ) );
BUF_X1 \keyboard/_1435_ ( .A(\keyboard/_0165_ ), .Z(\keyboard/_0336_ ) );
BUF_X1 \keyboard/_1436_ ( .A(\keyboard/_0189_ ), .Z(\keyboard/_0020_ ) );
BUF_X1 \keyboard/_1437_ ( .A(\keyboard/_0166_ ), .Z(\keyboard/_0337_ ) );
BUF_X1 \keyboard/_1438_ ( .A(\keyboard/_0190_ ), .Z(\keyboard/_0021_ ) );
BUF_X1 \keyboard/_1439_ ( .A(\keyboard/_0167_ ), .Z(\keyboard/_0338_ ) );
BUF_X1 \keyboard/_1440_ ( .A(\keyboard/_0169_ ), .Z(\keyboard/_0000_ ) );
BUF_X1 \keyboard/_1441_ ( .A(\keyboard/_0170_ ), .Z(\keyboard/_0001_ ) );
BUF_X1 \keyboard/_1442_ ( .A(\keyboard/_0171_ ), .Z(\keyboard/_0002_ ) );
BUF_X1 \keyboard/_1443_ ( .A(\keyboard/_0172_ ), .Z(\keyboard/_0003_ ) );
BUF_X1 \keyboard/_1444_ ( .A(\keyboard/_0173_ ), .Z(\keyboard/_0004_ ) );
BUF_X1 \keyboard/_1445_ ( .A(\keyboard/_0174_ ), .Z(\keyboard/_0005_ ) );
BUF_X1 \keyboard/_1446_ ( .A(\keyboard/_0175_ ), .Z(\keyboard/_0006_ ) );
BUF_X1 \keyboard/_1447_ ( .A(\keyboard/_0176_ ), .Z(\keyboard/_0007_ ) );
BUF_X1 \keyboard/_1448_ ( .A(\keyboard/_0177_ ), .Z(\keyboard/_0008_ ) );
BUF_X1 \keyboard/_1449_ ( .A(\keyboard/_0168_ ), .Z(\keyboard/_0339_ ) );
BUF_X1 \keyboard/_1450_ ( .A(\keyboard/_0178_ ), .Z(\keyboard/_0009_ ) );
DFF_X1 \keyboard/_1451_ ( .D(\keyboard/_0000_ ), .CK(clock ), .Q(\keyboard/buffer[0] ), .QN(\keyboard/_0167_ ) );
DFF_X1 \keyboard/_1452_ ( .D(\keyboard/_0001_ ), .CK(clock ), .Q(\keyboard/buffer[1] ), .QN(\keyboard/_0096_ ) );
DFF_X1 \keyboard/_1453_ ( .D(\keyboard/_0002_ ), .CK(clock ), .Q(\keyboard/buffer[2] ), .QN(\keyboard/_0098_ ) );
DFF_X1 \keyboard/_1454_ ( .D(\keyboard/_0003_ ), .CK(clock ), .Q(\keyboard/buffer[3] ), .QN(\keyboard/_0100_ ) );
DFF_X1 \keyboard/_1455_ ( .D(\keyboard/_0004_ ), .CK(clock ), .Q(\keyboard/buffer[4] ), .QN(\keyboard/_0102_ ) );
DFF_X1 \keyboard/_1456_ ( .D(\keyboard/_0005_ ), .CK(clock ), .Q(\keyboard/buffer[5] ), .QN(\keyboard/_0104_ ) );
DFF_X1 \keyboard/_1457_ ( .D(\keyboard/_0006_ ), .CK(clock ), .Q(\keyboard/buffer[6] ), .QN(\keyboard/_0106_ ) );
DFF_X1 \keyboard/_1458_ ( .D(\keyboard/_0007_ ), .CK(clock ), .Q(\keyboard/buffer[7] ), .QN(\keyboard/_0108_ ) );
DFF_X1 \keyboard/_1459_ ( .D(\keyboard/_0008_ ), .CK(clock ), .Q(\keyboard/buffer[8] ), .QN(\keyboard/_0110_ ) );
DFF_X1 \keyboard/_1460_ ( .D(\keyboard/_0009_ ), .CK(clock ), .Q(\keyboard/buffer[9] ), .QN(\keyboard/_0168_ ) );
DFF_X1 \keyboard/_1461_ ( .D(\keyboard/_0014_ ), .CK(clock ), .Q(\keyboard/fifo_0[0] ), .QN(\keyboard/_0159_ ) );
DFF_X1 \keyboard/_1462_ ( .D(\keyboard/_0015_ ), .CK(clock ), .Q(\keyboard/fifo_0[1] ), .QN(\keyboard/_0160_ ) );
DFF_X1 \keyboard/_1463_ ( .D(\keyboard/_0016_ ), .CK(clock ), .Q(\keyboard/fifo_0[2] ), .QN(\keyboard/_0161_ ) );
DFF_X1 \keyboard/_1464_ ( .D(\keyboard/_0017_ ), .CK(clock ), .Q(\keyboard/fifo_0[3] ), .QN(\keyboard/_0162_ ) );
DFF_X1 \keyboard/_1465_ ( .D(\keyboard/_0018_ ), .CK(clock ), .Q(\keyboard/fifo_0[4] ), .QN(\keyboard/_0163_ ) );
DFF_X1 \keyboard/_1466_ ( .D(\keyboard/_0019_ ), .CK(clock ), .Q(\keyboard/fifo_0[5] ), .QN(\keyboard/_0164_ ) );
DFF_X1 \keyboard/_1467_ ( .D(\keyboard/_0020_ ), .CK(clock ), .Q(\keyboard/fifo_0[6] ), .QN(\keyboard/_0165_ ) );
DFF_X1 \keyboard/_1468_ ( .D(\keyboard/_0021_ ), .CK(clock ), .Q(\keyboard/fifo_0[7] ), .QN(\keyboard/_0166_ ) );
DFF_X1 \keyboard/_1469_ ( .D(\keyboard/_0022_ ), .CK(clock ), .Q(\keyboard/fifo_1[0] ), .QN(\keyboard/_0151_ ) );
DFF_X1 \keyboard/_1470_ ( .D(\keyboard/_0023_ ), .CK(clock ), .Q(\keyboard/fifo_1[1] ), .QN(\keyboard/_0152_ ) );
DFF_X1 \keyboard/_1471_ ( .D(\keyboard/_0024_ ), .CK(clock ), .Q(\keyboard/fifo_1[2] ), .QN(\keyboard/_0153_ ) );
DFF_X1 \keyboard/_1472_ ( .D(\keyboard/_0025_ ), .CK(clock ), .Q(\keyboard/fifo_1[3] ), .QN(\keyboard/_0154_ ) );
DFF_X1 \keyboard/_1473_ ( .D(\keyboard/_0026_ ), .CK(clock ), .Q(\keyboard/fifo_1[4] ), .QN(\keyboard/_0155_ ) );
DFF_X1 \keyboard/_1474_ ( .D(\keyboard/_0027_ ), .CK(clock ), .Q(\keyboard/fifo_1[5] ), .QN(\keyboard/_0156_ ) );
DFF_X1 \keyboard/_1475_ ( .D(\keyboard/_0028_ ), .CK(clock ), .Q(\keyboard/fifo_1[6] ), .QN(\keyboard/_0157_ ) );
DFF_X1 \keyboard/_1476_ ( .D(\keyboard/_0029_ ), .CK(clock ), .Q(\keyboard/fifo_1[7] ), .QN(\keyboard/_0158_ ) );
DFF_X1 \keyboard/_1477_ ( .D(\keyboard/_0030_ ), .CK(clock ), .Q(\keyboard/fifo_2[0] ), .QN(\keyboard/_0143_ ) );
DFF_X1 \keyboard/_1478_ ( .D(\keyboard/_0031_ ), .CK(clock ), .Q(\keyboard/fifo_2[1] ), .QN(\keyboard/_0144_ ) );
DFF_X1 \keyboard/_1479_ ( .D(\keyboard/_0032_ ), .CK(clock ), .Q(\keyboard/fifo_2[2] ), .QN(\keyboard/_0145_ ) );
DFF_X1 \keyboard/_1480_ ( .D(\keyboard/_0033_ ), .CK(clock ), .Q(\keyboard/fifo_2[3] ), .QN(\keyboard/_0146_ ) );
DFF_X1 \keyboard/_1481_ ( .D(\keyboard/_0034_ ), .CK(clock ), .Q(\keyboard/fifo_2[4] ), .QN(\keyboard/_0147_ ) );
DFF_X1 \keyboard/_1482_ ( .D(\keyboard/_0035_ ), .CK(clock ), .Q(\keyboard/fifo_2[5] ), .QN(\keyboard/_0148_ ) );
DFF_X1 \keyboard/_1483_ ( .D(\keyboard/_0036_ ), .CK(clock ), .Q(\keyboard/fifo_2[6] ), .QN(\keyboard/_0149_ ) );
DFF_X1 \keyboard/_1484_ ( .D(\keyboard/_0037_ ), .CK(clock ), .Q(\keyboard/fifo_2[7] ), .QN(\keyboard/_0150_ ) );
DFF_X1 \keyboard/_1485_ ( .D(\keyboard/_0038_ ), .CK(clock ), .Q(\keyboard/fifo_3[0] ), .QN(\keyboard/_0135_ ) );
DFF_X1 \keyboard/_1486_ ( .D(\keyboard/_0039_ ), .CK(clock ), .Q(\keyboard/fifo_3[1] ), .QN(\keyboard/_0136_ ) );
DFF_X1 \keyboard/_1487_ ( .D(\keyboard/_0040_ ), .CK(clock ), .Q(\keyboard/fifo_3[2] ), .QN(\keyboard/_0137_ ) );
DFF_X1 \keyboard/_1488_ ( .D(\keyboard/_0041_ ), .CK(clock ), .Q(\keyboard/fifo_3[3] ), .QN(\keyboard/_0138_ ) );
DFF_X1 \keyboard/_1489_ ( .D(\keyboard/_0042_ ), .CK(clock ), .Q(\keyboard/fifo_3[4] ), .QN(\keyboard/_0139_ ) );
DFF_X1 \keyboard/_1490_ ( .D(\keyboard/_0043_ ), .CK(clock ), .Q(\keyboard/fifo_3[5] ), .QN(\keyboard/_0140_ ) );
DFF_X1 \keyboard/_1491_ ( .D(\keyboard/_0044_ ), .CK(clock ), .Q(\keyboard/fifo_3[6] ), .QN(\keyboard/_0141_ ) );
DFF_X1 \keyboard/_1492_ ( .D(\keyboard/_0045_ ), .CK(clock ), .Q(\keyboard/fifo_3[7] ), .QN(\keyboard/_0142_ ) );
DFF_X1 \keyboard/_1493_ ( .D(\keyboard/_0046_ ), .CK(clock ), .Q(\keyboard/fifo_4[0] ), .QN(\keyboard/_0127_ ) );
DFF_X1 \keyboard/_1494_ ( .D(\keyboard/_0047_ ), .CK(clock ), .Q(\keyboard/fifo_4[1] ), .QN(\keyboard/_0128_ ) );
DFF_X1 \keyboard/_1495_ ( .D(\keyboard/_0048_ ), .CK(clock ), .Q(\keyboard/fifo_4[2] ), .QN(\keyboard/_0129_ ) );
DFF_X1 \keyboard/_1496_ ( .D(\keyboard/_0049_ ), .CK(clock ), .Q(\keyboard/fifo_4[3] ), .QN(\keyboard/_0130_ ) );
DFF_X1 \keyboard/_1497_ ( .D(\keyboard/_0050_ ), .CK(clock ), .Q(\keyboard/fifo_4[4] ), .QN(\keyboard/_0131_ ) );
DFF_X1 \keyboard/_1498_ ( .D(\keyboard/_0051_ ), .CK(clock ), .Q(\keyboard/fifo_4[5] ), .QN(\keyboard/_0132_ ) );
DFF_X1 \keyboard/_1499_ ( .D(\keyboard/_0052_ ), .CK(clock ), .Q(\keyboard/fifo_4[6] ), .QN(\keyboard/_0133_ ) );
DFF_X1 \keyboard/_1500_ ( .D(\keyboard/_0053_ ), .CK(clock ), .Q(\keyboard/fifo_4[7] ), .QN(\keyboard/_0134_ ) );
DFF_X1 \keyboard/_1501_ ( .D(\keyboard/_0054_ ), .CK(clock ), .Q(\keyboard/fifo_5[0] ), .QN(\keyboard/_0119_ ) );
DFF_X1 \keyboard/_1502_ ( .D(\keyboard/_0055_ ), .CK(clock ), .Q(\keyboard/fifo_5[1] ), .QN(\keyboard/_0120_ ) );
DFF_X1 \keyboard/_1503_ ( .D(\keyboard/_0056_ ), .CK(clock ), .Q(\keyboard/fifo_5[2] ), .QN(\keyboard/_0121_ ) );
DFF_X1 \keyboard/_1504_ ( .D(\keyboard/_0057_ ), .CK(clock ), .Q(\keyboard/fifo_5[3] ), .QN(\keyboard/_0122_ ) );
DFF_X1 \keyboard/_1505_ ( .D(\keyboard/_0058_ ), .CK(clock ), .Q(\keyboard/fifo_5[4] ), .QN(\keyboard/_0123_ ) );
DFF_X1 \keyboard/_1506_ ( .D(\keyboard/_0059_ ), .CK(clock ), .Q(\keyboard/fifo_5[5] ), .QN(\keyboard/_0124_ ) );
DFF_X1 \keyboard/_1507_ ( .D(\keyboard/_0060_ ), .CK(clock ), .Q(\keyboard/fifo_5[6] ), .QN(\keyboard/_0125_ ) );
DFF_X1 \keyboard/_1508_ ( .D(\keyboard/_0061_ ), .CK(clock ), .Q(\keyboard/fifo_5[7] ), .QN(\keyboard/_0126_ ) );
DFF_X1 \keyboard/_1509_ ( .D(\keyboard/_0062_ ), .CK(clock ), .Q(\keyboard/fifo_6[0] ), .QN(\keyboard/_0111_ ) );
DFF_X1 \keyboard/_1510_ ( .D(\keyboard/_0063_ ), .CK(clock ), .Q(\keyboard/fifo_6[1] ), .QN(\keyboard/_0112_ ) );
DFF_X1 \keyboard/_1511_ ( .D(\keyboard/_0064_ ), .CK(clock ), .Q(\keyboard/fifo_6[2] ), .QN(\keyboard/_0113_ ) );
DFF_X1 \keyboard/_1512_ ( .D(\keyboard/_0065_ ), .CK(clock ), .Q(\keyboard/fifo_6[3] ), .QN(\keyboard/_0114_ ) );
DFF_X1 \keyboard/_1513_ ( .D(\keyboard/_0066_ ), .CK(clock ), .Q(\keyboard/fifo_6[4] ), .QN(\keyboard/_0115_ ) );
DFF_X1 \keyboard/_1514_ ( .D(\keyboard/_0067_ ), .CK(clock ), .Q(\keyboard/fifo_6[5] ), .QN(\keyboard/_0116_ ) );
DFF_X1 \keyboard/_1515_ ( .D(\keyboard/_0068_ ), .CK(clock ), .Q(\keyboard/fifo_6[6] ), .QN(\keyboard/_0117_ ) );
DFF_X1 \keyboard/_1516_ ( .D(\keyboard/_0069_ ), .CK(clock ), .Q(\keyboard/fifo_6[7] ), .QN(\keyboard/_0118_ ) );
DFF_X1 \keyboard/_1517_ ( .D(\keyboard/_0070_ ), .CK(clock ), .Q(\keyboard/fifo_7[0] ), .QN(\keyboard/_0095_ ) );
DFF_X1 \keyboard/_1518_ ( .D(\keyboard/_0071_ ), .CK(clock ), .Q(\keyboard/fifo_7[1] ), .QN(\keyboard/_0097_ ) );
DFF_X1 \keyboard/_1519_ ( .D(\keyboard/_0072_ ), .CK(clock ), .Q(\keyboard/fifo_7[2] ), .QN(\keyboard/_0099_ ) );
DFF_X1 \keyboard/_1520_ ( .D(\keyboard/_0073_ ), .CK(clock ), .Q(\keyboard/fifo_7[3] ), .QN(\keyboard/_0101_ ) );
DFF_X1 \keyboard/_1521_ ( .D(\keyboard/_0074_ ), .CK(clock ), .Q(\keyboard/fifo_7[4] ), .QN(\keyboard/_0103_ ) );
DFF_X1 \keyboard/_1522_ ( .D(\keyboard/_0075_ ), .CK(clock ), .Q(\keyboard/fifo_7[5] ), .QN(\keyboard/_0105_ ) );
DFF_X1 \keyboard/_1523_ ( .D(\keyboard/_0076_ ), .CK(clock ), .Q(\keyboard/fifo_7[6] ), .QN(\keyboard/_0107_ ) );
DFF_X1 \keyboard/_1524_ ( .D(\keyboard/_0077_ ), .CK(clock ), .Q(\keyboard/fifo_7[7] ), .QN(\keyboard/_0109_ ) );
DFF_X1 \keyboard/_1525_ ( .D(\keyboard/_0085_ ), .CK(clock ), .Q(\keyboard/w_ptr[0] ), .QN(\keyboard/_0094_ ) );
DFF_X1 \keyboard/_1526_ ( .D(\keyboard/_0086_ ), .CK(clock ), .Q(\keyboard/w_ptr[1] ), .QN(\keyboard/_0089_ ) );
DFF_X1 \keyboard/_1527_ ( .D(\keyboard/_0087_ ), .CK(clock ), .Q(\keyboard/w_ptr[2] ), .QN(\keyboard/_0090_ ) );
DFF_X1 \keyboard/_1528_ ( .D(\keyboard/_0081_ ), .CK(clock ), .Q(\keyboard/r_ptr[0] ), .QN(\keyboard/_0757_ ) );
DFF_X1 \keyboard/_1529_ ( .D(\keyboard/_0082_ ), .CK(clock ), .Q(\keyboard/r_ptr[1] ), .QN(\keyboard/_0093_ ) );
DFF_X1 \keyboard/_1530_ ( .D(\keyboard/_0083_ ), .CK(clock ), .Q(\keyboard/r_ptr[2] ), .QN(\keyboard/_0088_ ) );
DFF_X1 \keyboard/_1531_ ( .D(\keyboard/_0010_ ), .CK(clock ), .Q(\keyboard/count[0] ), .QN(\keyboard/_0091_ ) );
DFF_X1 \keyboard/_1532_ ( .D(\keyboard/_0011_ ), .CK(clock ), .Q(\keyboard/count[1] ), .QN(\keyboard/_0758_ ) );
DFF_X1 \keyboard/_1533_ ( .D(\keyboard/_0012_ ), .CK(clock ), .Q(\keyboard/count[2] ), .QN(\keyboard/_0759_ ) );
DFF_X1 \keyboard/_1534_ ( .D(\keyboard/_0013_ ), .CK(clock ), .Q(\keyboard/count[3] ), .QN(\keyboard/_0092_ ) );
DFF_X1 \keyboard/_1535_ ( .D(\keyboard/_0084_ ), .CK(clock ), .Q(keyboard_io_ready ), .QN(\keyboard/_0760_ ) );
DFF_X1 \keyboard/_1536_ ( .D(\keyboard/_0078_ ), .CK(clock ), .Q(\keyboard/_ps2_clk_sync_T_1[1] ), .QN(\keyboard/_0761_ ) );
DFF_X1 \keyboard/_1537_ ( .D(\keyboard/_0079_ ), .CK(clock ), .Q(\keyboard/_ps2_clk_sync_T_1[2] ), .QN(\keyboard/_0762_ ) );
DFF_X1 \keyboard/_1538_ ( .D(\keyboard/_0080_ ), .CK(clock ), .Q(\keyboard/ps2_clk_sync[2] ), .QN(\keyboard/_0763_ ) );
INV_X32 \seg0/_062_ ( .A(\seg0/_003_ ), .ZN(\seg0/_013_ ) );
NOR2_X4 \seg0/_063_ ( .A1(\seg0/_013_ ), .A2(\seg0/_005_ ), .ZN(\seg0/_014_ ) );
AND2_X4 \seg0/_064_ ( .A1(\seg0/_014_ ), .A2(\seg0/_004_ ), .ZN(\seg0/_015_ ) );
INV_X32 \seg0/_065_ ( .A(\seg0/_001_ ), .ZN(\seg0/_016_ ) );
NOR2_X4 \seg0/_066_ ( .A1(\seg0/_016_ ), .A2(\seg0/_002_ ), .ZN(\seg0/_017_ ) );
AND2_X2 \seg0/_067_ ( .A1(\seg0/_015_ ), .A2(\seg0/_017_ ), .ZN(\seg0/_018_ ) );
NOR2_X4 \seg0/_068_ ( .A1(\seg0/_005_ ), .A2(\seg0/_003_ ), .ZN(\seg0/_019_ ) );
AND2_X1 \seg0/_069_ ( .A1(\seg0/_019_ ), .A2(\seg0/_004_ ), .ZN(\seg0/_020_ ) );
NOR2_X2 \seg0/_070_ ( .A1(\seg0/_018_ ), .A2(\seg0/_020_ ), .ZN(\seg0/_021_ ) );
AND2_X4 \seg0/_071_ ( .A1(\seg0/_002_ ), .A2(\seg0/_001_ ), .ZN(\seg0/_022_ ) );
INV_X4 \seg0/_072_ ( .A(\seg0/_022_ ), .ZN(\seg0/_023_ ) );
INV_X32 \seg0/_073_ ( .A(\seg0/_004_ ), .ZN(\seg0/_024_ ) );
NAND3_X1 \seg0/_074_ ( .A1(\seg0/_023_ ), .A2(\seg0/_024_ ), .A3(\seg0/_014_ ), .ZN(\seg0/_025_ ) );
AND2_X4 \seg0/_075_ ( .A1(\seg0/_019_ ), .A2(\seg0/_024_ ), .ZN(\seg0/_026_ ) );
NAND2_X1 \seg0/_076_ ( .A1(\seg0/_026_ ), .A2(\seg0/_022_ ), .ZN(\seg0/_027_ ) );
NAND2_X1 \seg0/_077_ ( .A1(\seg0/_015_ ), .A2(\seg0/_002_ ), .ZN(\seg0/_028_ ) );
NAND4_X1 \seg0/_078_ ( .A1(\seg0/_021_ ), .A2(\seg0/_025_ ), .A3(\seg0/_027_ ), .A4(\seg0/_028_ ), .ZN(\seg0/_029_ ) );
INV_X16 \seg0/_079_ ( .A(\seg0/_002_ ), .ZN(\seg0/_030_ ) );
NOR2_X4 \seg0/_080_ ( .A1(\seg0/_030_ ), .A2(\seg0/_001_ ), .ZN(\seg0/_031_ ) );
AND2_X4 \seg0/_081_ ( .A1(\seg0/_026_ ), .A2(\seg0/_031_ ), .ZN(\seg0/_032_ ) );
OAI21_X1 \seg0/_082_ ( .A(\seg0/_000_ ), .B1(\seg0/_029_ ), .B2(\seg0/_032_ ), .ZN(\seg0/_006_ ) );
INV_X1 \seg0/_083_ ( .A(\seg0/_017_ ), .ZN(\seg0/_033_ ) );
AND2_X4 \seg0/_084_ ( .A1(\seg0/_015_ ), .A2(\seg0/_033_ ), .ZN(\seg0/_034_ ) );
AND3_X2 \seg0/_085_ ( .A1(\seg0/_023_ ), .A2(\seg0/_004_ ), .A3(\seg0/_019_ ), .ZN(\seg0/_035_ ) );
NOR2_X2 \seg0/_086_ ( .A1(\seg0/_034_ ), .A2(\seg0/_035_ ), .ZN(\seg0/_036_ ) );
NAND2_X1 \seg0/_087_ ( .A1(\seg0/_020_ ), .A2(\seg0/_022_ ), .ZN(\seg0/_037_ ) );
NOR2_X4 \seg0/_088_ ( .A1(\seg0/_002_ ), .A2(\seg0/_001_ ), .ZN(\seg0/_038_ ) );
NAND2_X1 \seg0/_089_ ( .A1(\seg0/_026_ ), .A2(\seg0/_038_ ), .ZN(\seg0/_039_ ) );
NAND4_X1 \seg0/_090_ ( .A1(\seg0/_036_ ), .A2(\seg0/_037_ ), .A3(\seg0/_025_ ), .A4(\seg0/_039_ ), .ZN(\seg0/_040_ ) );
NAND2_X1 \seg0/_091_ ( .A1(\seg0/_040_ ), .A2(\seg0/_000_ ), .ZN(\seg0/_007_ ) );
AND2_X1 \seg0/_092_ ( .A1(\seg0/_019_ ), .A2(\seg0/_038_ ), .ZN(\seg0/_041_ ) );
OR4_X4 \seg0/_093_ ( .A1(\seg0/_018_ ), .A2(\seg0/_034_ ), .A3(\seg0/_041_ ), .A4(\seg0/_032_ ), .ZN(\seg0/_042_ ) );
AND2_X1 \seg0/_094_ ( .A1(\seg0/_014_ ), .A2(\seg0/_024_ ), .ZN(\seg0/_043_ ) );
NAND2_X1 \seg0/_095_ ( .A1(\seg0/_043_ ), .A2(\seg0/_031_ ), .ZN(\seg0/_044_ ) );
NAND2_X1 \seg0/_096_ ( .A1(\seg0/_020_ ), .A2(\seg0/_031_ ), .ZN(\seg0/_045_ ) );
NAND3_X1 \seg0/_097_ ( .A1(\seg0/_044_ ), .A2(\seg0/_045_ ), .A3(\seg0/_037_ ), .ZN(\seg0/_046_ ) );
OAI21_X1 \seg0/_098_ ( .A(\seg0/_000_ ), .B1(\seg0/_042_ ), .B2(\seg0/_046_ ), .ZN(\seg0/_008_ ) );
INV_X1 \seg0/_099_ ( .A(\seg0/_043_ ), .ZN(\seg0/_047_ ) );
OAI21_X1 \seg0/_100_ ( .A(\seg0/_044_ ), .B1(\seg0/_047_ ), .B2(\seg0/_033_ ), .ZN(\seg0/_048_ ) );
NAND2_X1 \seg0/_101_ ( .A1(\seg0/_041_ ), .A2(\seg0/_004_ ), .ZN(\seg0/_049_ ) );
NAND2_X1 \seg0/_102_ ( .A1(\seg0/_026_ ), .A2(\seg0/_033_ ), .ZN(\seg0/_050_ ) );
NAND3_X1 \seg0/_103_ ( .A1(\seg0/_023_ ), .A2(\seg0/_004_ ), .A3(\seg0/_014_ ), .ZN(\seg0/_051_ ) );
NAND3_X1 \seg0/_104_ ( .A1(\seg0/_019_ ), .A2(\seg0/_001_ ), .A3(\seg0/_004_ ), .ZN(\seg0/_052_ ) );
NAND4_X1 \seg0/_105_ ( .A1(\seg0/_049_ ), .A2(\seg0/_050_ ), .A3(\seg0/_051_ ), .A4(\seg0/_052_ ), .ZN(\seg0/_053_ ) );
OAI21_X1 \seg0/_106_ ( .A(\seg0/_000_ ), .B1(\seg0/_048_ ), .B2(\seg0/_053_ ), .ZN(\seg0/_009_ ) );
INV_X1 \seg0/_107_ ( .A(\seg0/_021_ ), .ZN(\seg0/_054_ ) );
AOI211_X4 \seg0/_108_ ( .A(\seg0/_005_ ), .B(\seg0/_004_ ), .C1(\seg0/_031_ ), .C2(\seg0/_013_ ), .ZN(\seg0/_055_ ) );
OAI21_X1 \seg0/_109_ ( .A(\seg0/_000_ ), .B1(\seg0/_054_ ), .B2(\seg0/_055_ ), .ZN(\seg0/_010_ ) );
NAND3_X1 \seg0/_110_ ( .A1(\seg0/_014_ ), .A2(\seg0/_030_ ), .A3(\seg0/_024_ ), .ZN(\seg0/_056_ ) );
NOR2_X1 \seg0/_111_ ( .A1(\seg0/_056_ ), .A2(\seg0/_001_ ), .ZN(\seg0/_057_ ) );
OR3_X2 \seg0/_112_ ( .A1(\seg0/_018_ ), .A2(\seg0/_057_ ), .A3(\seg0/_035_ ), .ZN(\seg0/_058_ ) );
AOI211_X4 \seg0/_113_ ( .A(\seg0/_005_ ), .B(\seg0/_004_ ), .C1(\seg0/_023_ ), .C2(\seg0/_003_ ), .ZN(\seg0/_059_ ) );
OAI21_X1 \seg0/_114_ ( .A(\seg0/_000_ ), .B1(\seg0/_058_ ), .B2(\seg0/_059_ ), .ZN(\seg0/_011_ ) );
OAI211_X2 \seg0/_115_ ( .A(\seg0/_036_ ), .B(\seg0/_050_ ), .C1(\seg0/_038_ ), .C2(\seg0/_047_ ), .ZN(\seg0/_060_ ) );
NAND2_X1 \seg0/_116_ ( .A1(\seg0/_060_ ), .A2(\seg0/_000_ ), .ZN(\seg0/_012_ ) );
LOGIC1_X1 \seg0/_117_ ( .Z(\seg0/_061_ ) );
BUF_X1 \seg0/_118_ ( .A(\seg0/_061_ ), .Z(\io_seg_out_0[0] ) );
BUF_X1 \seg0/_119_ ( .A(display_en ), .Z(\seg0/_000_ ) );
BUF_X1 \seg0/_120_ ( .A(_194_ ), .Z(\seg0/_005_ ) );
BUF_X1 \seg0/_121_ ( .A(\seg0_in[1] ), .Z(\seg0/_002_ ) );
BUF_X1 \seg0/_122_ ( .A(\seg0_in[0] ), .Z(\seg0/_001_ ) );
BUF_X1 \seg0/_123_ ( .A(\seg0_in[3] ), .Z(\seg0/_004_ ) );
BUF_X1 \seg0/_124_ ( .A(\seg0_in[2] ), .Z(\seg0/_003_ ) );
BUF_X1 \seg0/_125_ ( .A(\seg0/_006_ ), .Z(\io_seg_out_0[1] ) );
BUF_X1 \seg0/_126_ ( .A(\seg0/_007_ ), .Z(\io_seg_out_0[2] ) );
BUF_X1 \seg0/_127_ ( .A(\seg0/_008_ ), .Z(\io_seg_out_0[3] ) );
BUF_X1 \seg0/_128_ ( .A(\seg0/_009_ ), .Z(\io_seg_out_0[4] ) );
BUF_X1 \seg0/_129_ ( .A(\seg0/_010_ ), .Z(\io_seg_out_0[5] ) );
BUF_X1 \seg0/_130_ ( .A(\seg0/_011_ ), .Z(\io_seg_out_0[6] ) );
BUF_X1 \seg0/_131_ ( .A(\seg0/_012_ ), .Z(\io_seg_out_0[7] ) );
INV_X32 \seg1/_062_ ( .A(\seg1/_003_ ), .ZN(\seg1/_013_ ) );
NOR2_X4 \seg1/_063_ ( .A1(\seg1/_013_ ), .A2(\seg1/_005_ ), .ZN(\seg1/_014_ ) );
AND2_X4 \seg1/_064_ ( .A1(\seg1/_014_ ), .A2(\seg1/_004_ ), .ZN(\seg1/_015_ ) );
INV_X32 \seg1/_065_ ( .A(\seg1/_001_ ), .ZN(\seg1/_016_ ) );
NOR2_X4 \seg1/_066_ ( .A1(\seg1/_016_ ), .A2(\seg1/_002_ ), .ZN(\seg1/_017_ ) );
AND2_X2 \seg1/_067_ ( .A1(\seg1/_015_ ), .A2(\seg1/_017_ ), .ZN(\seg1/_018_ ) );
NOR2_X4 \seg1/_068_ ( .A1(\seg1/_005_ ), .A2(\seg1/_003_ ), .ZN(\seg1/_019_ ) );
AND2_X1 \seg1/_069_ ( .A1(\seg1/_019_ ), .A2(\seg1/_004_ ), .ZN(\seg1/_020_ ) );
NOR2_X2 \seg1/_070_ ( .A1(\seg1/_018_ ), .A2(\seg1/_020_ ), .ZN(\seg1/_021_ ) );
AND2_X4 \seg1/_071_ ( .A1(\seg1/_002_ ), .A2(\seg1/_001_ ), .ZN(\seg1/_022_ ) );
INV_X4 \seg1/_072_ ( .A(\seg1/_022_ ), .ZN(\seg1/_023_ ) );
INV_X32 \seg1/_073_ ( .A(\seg1/_004_ ), .ZN(\seg1/_024_ ) );
NAND3_X1 \seg1/_074_ ( .A1(\seg1/_023_ ), .A2(\seg1/_024_ ), .A3(\seg1/_014_ ), .ZN(\seg1/_025_ ) );
AND2_X4 \seg1/_075_ ( .A1(\seg1/_019_ ), .A2(\seg1/_024_ ), .ZN(\seg1/_026_ ) );
NAND2_X1 \seg1/_076_ ( .A1(\seg1/_026_ ), .A2(\seg1/_022_ ), .ZN(\seg1/_027_ ) );
NAND2_X1 \seg1/_077_ ( .A1(\seg1/_015_ ), .A2(\seg1/_002_ ), .ZN(\seg1/_028_ ) );
NAND4_X1 \seg1/_078_ ( .A1(\seg1/_021_ ), .A2(\seg1/_025_ ), .A3(\seg1/_027_ ), .A4(\seg1/_028_ ), .ZN(\seg1/_029_ ) );
INV_X16 \seg1/_079_ ( .A(\seg1/_002_ ), .ZN(\seg1/_030_ ) );
NOR2_X4 \seg1/_080_ ( .A1(\seg1/_030_ ), .A2(\seg1/_001_ ), .ZN(\seg1/_031_ ) );
AND2_X4 \seg1/_081_ ( .A1(\seg1/_026_ ), .A2(\seg1/_031_ ), .ZN(\seg1/_032_ ) );
OAI21_X1 \seg1/_082_ ( .A(\seg1/_000_ ), .B1(\seg1/_029_ ), .B2(\seg1/_032_ ), .ZN(\seg1/_006_ ) );
INV_X1 \seg1/_083_ ( .A(\seg1/_017_ ), .ZN(\seg1/_033_ ) );
AND2_X4 \seg1/_084_ ( .A1(\seg1/_015_ ), .A2(\seg1/_033_ ), .ZN(\seg1/_034_ ) );
AND3_X2 \seg1/_085_ ( .A1(\seg1/_023_ ), .A2(\seg1/_004_ ), .A3(\seg1/_019_ ), .ZN(\seg1/_035_ ) );
NOR2_X2 \seg1/_086_ ( .A1(\seg1/_034_ ), .A2(\seg1/_035_ ), .ZN(\seg1/_036_ ) );
NAND2_X1 \seg1/_087_ ( .A1(\seg1/_020_ ), .A2(\seg1/_022_ ), .ZN(\seg1/_037_ ) );
NOR2_X4 \seg1/_088_ ( .A1(\seg1/_002_ ), .A2(\seg1/_001_ ), .ZN(\seg1/_038_ ) );
NAND2_X1 \seg1/_089_ ( .A1(\seg1/_026_ ), .A2(\seg1/_038_ ), .ZN(\seg1/_039_ ) );
NAND4_X1 \seg1/_090_ ( .A1(\seg1/_036_ ), .A2(\seg1/_037_ ), .A3(\seg1/_025_ ), .A4(\seg1/_039_ ), .ZN(\seg1/_040_ ) );
NAND2_X1 \seg1/_091_ ( .A1(\seg1/_040_ ), .A2(\seg1/_000_ ), .ZN(\seg1/_007_ ) );
AND2_X1 \seg1/_092_ ( .A1(\seg1/_019_ ), .A2(\seg1/_038_ ), .ZN(\seg1/_041_ ) );
OR4_X4 \seg1/_093_ ( .A1(\seg1/_018_ ), .A2(\seg1/_034_ ), .A3(\seg1/_041_ ), .A4(\seg1/_032_ ), .ZN(\seg1/_042_ ) );
AND2_X1 \seg1/_094_ ( .A1(\seg1/_014_ ), .A2(\seg1/_024_ ), .ZN(\seg1/_043_ ) );
NAND2_X1 \seg1/_095_ ( .A1(\seg1/_043_ ), .A2(\seg1/_031_ ), .ZN(\seg1/_044_ ) );
NAND2_X1 \seg1/_096_ ( .A1(\seg1/_020_ ), .A2(\seg1/_031_ ), .ZN(\seg1/_045_ ) );
NAND3_X1 \seg1/_097_ ( .A1(\seg1/_044_ ), .A2(\seg1/_045_ ), .A3(\seg1/_037_ ), .ZN(\seg1/_046_ ) );
OAI21_X1 \seg1/_098_ ( .A(\seg1/_000_ ), .B1(\seg1/_042_ ), .B2(\seg1/_046_ ), .ZN(\seg1/_008_ ) );
INV_X1 \seg1/_099_ ( .A(\seg1/_043_ ), .ZN(\seg1/_047_ ) );
OAI21_X1 \seg1/_100_ ( .A(\seg1/_044_ ), .B1(\seg1/_047_ ), .B2(\seg1/_033_ ), .ZN(\seg1/_048_ ) );
NAND2_X1 \seg1/_101_ ( .A1(\seg1/_041_ ), .A2(\seg1/_004_ ), .ZN(\seg1/_049_ ) );
NAND2_X1 \seg1/_102_ ( .A1(\seg1/_026_ ), .A2(\seg1/_033_ ), .ZN(\seg1/_050_ ) );
NAND3_X1 \seg1/_103_ ( .A1(\seg1/_023_ ), .A2(\seg1/_004_ ), .A3(\seg1/_014_ ), .ZN(\seg1/_051_ ) );
NAND3_X1 \seg1/_104_ ( .A1(\seg1/_019_ ), .A2(\seg1/_001_ ), .A3(\seg1/_004_ ), .ZN(\seg1/_052_ ) );
NAND4_X1 \seg1/_105_ ( .A1(\seg1/_049_ ), .A2(\seg1/_050_ ), .A3(\seg1/_051_ ), .A4(\seg1/_052_ ), .ZN(\seg1/_053_ ) );
OAI21_X1 \seg1/_106_ ( .A(\seg1/_000_ ), .B1(\seg1/_048_ ), .B2(\seg1/_053_ ), .ZN(\seg1/_009_ ) );
INV_X1 \seg1/_107_ ( .A(\seg1/_021_ ), .ZN(\seg1/_054_ ) );
AOI211_X4 \seg1/_108_ ( .A(\seg1/_005_ ), .B(\seg1/_004_ ), .C1(\seg1/_031_ ), .C2(\seg1/_013_ ), .ZN(\seg1/_055_ ) );
OAI21_X1 \seg1/_109_ ( .A(\seg1/_000_ ), .B1(\seg1/_054_ ), .B2(\seg1/_055_ ), .ZN(\seg1/_010_ ) );
NAND3_X1 \seg1/_110_ ( .A1(\seg1/_014_ ), .A2(\seg1/_030_ ), .A3(\seg1/_024_ ), .ZN(\seg1/_056_ ) );
NOR2_X1 \seg1/_111_ ( .A1(\seg1/_056_ ), .A2(\seg1/_001_ ), .ZN(\seg1/_057_ ) );
OR3_X2 \seg1/_112_ ( .A1(\seg1/_018_ ), .A2(\seg1/_057_ ), .A3(\seg1/_035_ ), .ZN(\seg1/_058_ ) );
AOI211_X4 \seg1/_113_ ( .A(\seg1/_005_ ), .B(\seg1/_004_ ), .C1(\seg1/_023_ ), .C2(\seg1/_003_ ), .ZN(\seg1/_059_ ) );
OAI21_X1 \seg1/_114_ ( .A(\seg1/_000_ ), .B1(\seg1/_058_ ), .B2(\seg1/_059_ ), .ZN(\seg1/_011_ ) );
OAI211_X2 \seg1/_115_ ( .A(\seg1/_036_ ), .B(\seg1/_050_ ), .C1(\seg1/_038_ ), .C2(\seg1/_047_ ), .ZN(\seg1/_060_ ) );
NAND2_X1 \seg1/_116_ ( .A1(\seg1/_060_ ), .A2(\seg1/_000_ ), .ZN(\seg1/_012_ ) );
LOGIC1_X1 \seg1/_117_ ( .Z(\seg1/_061_ ) );
BUF_X1 \seg1/_118_ ( .A(\seg1/_061_ ), .Z(\io_seg_out_1[0] ) );
BUF_X1 \seg1/_119_ ( .A(display_en ), .Z(\seg1/_000_ ) );
BUF_X1 \seg1/_120_ ( .A(_194_ ), .Z(\seg1/_005_ ) );
BUF_X1 \seg1/_121_ ( .A(\seg1_in[1] ), .Z(\seg1/_002_ ) );
BUF_X1 \seg1/_122_ ( .A(\seg1_in[0] ), .Z(\seg1/_001_ ) );
BUF_X1 \seg1/_123_ ( .A(\seg1_in[3] ), .Z(\seg1/_004_ ) );
BUF_X1 \seg1/_124_ ( .A(\seg1_in[2] ), .Z(\seg1/_003_ ) );
BUF_X1 \seg1/_125_ ( .A(\seg1/_006_ ), .Z(\io_seg_out_1[1] ) );
BUF_X1 \seg1/_126_ ( .A(\seg1/_007_ ), .Z(\io_seg_out_1[2] ) );
BUF_X1 \seg1/_127_ ( .A(\seg1/_008_ ), .Z(\io_seg_out_1[3] ) );
BUF_X1 \seg1/_128_ ( .A(\seg1/_009_ ), .Z(\io_seg_out_1[4] ) );
BUF_X1 \seg1/_129_ ( .A(\seg1/_010_ ), .Z(\io_seg_out_1[5] ) );
BUF_X1 \seg1/_130_ ( .A(\seg1/_011_ ), .Z(\io_seg_out_1[6] ) );
BUF_X1 \seg1/_131_ ( .A(\seg1/_012_ ), .Z(\io_seg_out_1[7] ) );
INV_X32 \seg2/_062_ ( .A(\seg2/_003_ ), .ZN(\seg2/_013_ ) );
NOR2_X4 \seg2/_063_ ( .A1(\seg2/_013_ ), .A2(\seg2/_005_ ), .ZN(\seg2/_014_ ) );
AND2_X4 \seg2/_064_ ( .A1(\seg2/_014_ ), .A2(\seg2/_004_ ), .ZN(\seg2/_015_ ) );
INV_X32 \seg2/_065_ ( .A(\seg2/_001_ ), .ZN(\seg2/_016_ ) );
NOR2_X4 \seg2/_066_ ( .A1(\seg2/_016_ ), .A2(\seg2/_002_ ), .ZN(\seg2/_017_ ) );
AND2_X2 \seg2/_067_ ( .A1(\seg2/_015_ ), .A2(\seg2/_017_ ), .ZN(\seg2/_018_ ) );
NOR2_X4 \seg2/_068_ ( .A1(\seg2/_005_ ), .A2(\seg2/_003_ ), .ZN(\seg2/_019_ ) );
AND2_X1 \seg2/_069_ ( .A1(\seg2/_019_ ), .A2(\seg2/_004_ ), .ZN(\seg2/_020_ ) );
NOR2_X2 \seg2/_070_ ( .A1(\seg2/_018_ ), .A2(\seg2/_020_ ), .ZN(\seg2/_021_ ) );
AND2_X4 \seg2/_071_ ( .A1(\seg2/_002_ ), .A2(\seg2/_001_ ), .ZN(\seg2/_022_ ) );
INV_X4 \seg2/_072_ ( .A(\seg2/_022_ ), .ZN(\seg2/_023_ ) );
INV_X32 \seg2/_073_ ( .A(\seg2/_004_ ), .ZN(\seg2/_024_ ) );
NAND3_X1 \seg2/_074_ ( .A1(\seg2/_023_ ), .A2(\seg2/_024_ ), .A3(\seg2/_014_ ), .ZN(\seg2/_025_ ) );
AND2_X4 \seg2/_075_ ( .A1(\seg2/_019_ ), .A2(\seg2/_024_ ), .ZN(\seg2/_026_ ) );
NAND2_X1 \seg2/_076_ ( .A1(\seg2/_026_ ), .A2(\seg2/_022_ ), .ZN(\seg2/_027_ ) );
NAND2_X1 \seg2/_077_ ( .A1(\seg2/_015_ ), .A2(\seg2/_002_ ), .ZN(\seg2/_028_ ) );
NAND4_X1 \seg2/_078_ ( .A1(\seg2/_021_ ), .A2(\seg2/_025_ ), .A3(\seg2/_027_ ), .A4(\seg2/_028_ ), .ZN(\seg2/_029_ ) );
INV_X16 \seg2/_079_ ( .A(\seg2/_002_ ), .ZN(\seg2/_030_ ) );
NOR2_X4 \seg2/_080_ ( .A1(\seg2/_030_ ), .A2(\seg2/_001_ ), .ZN(\seg2/_031_ ) );
AND2_X4 \seg2/_081_ ( .A1(\seg2/_026_ ), .A2(\seg2/_031_ ), .ZN(\seg2/_032_ ) );
OAI21_X1 \seg2/_082_ ( .A(\seg2/_000_ ), .B1(\seg2/_029_ ), .B2(\seg2/_032_ ), .ZN(\seg2/_006_ ) );
INV_X1 \seg2/_083_ ( .A(\seg2/_017_ ), .ZN(\seg2/_033_ ) );
AND2_X4 \seg2/_084_ ( .A1(\seg2/_015_ ), .A2(\seg2/_033_ ), .ZN(\seg2/_034_ ) );
AND3_X2 \seg2/_085_ ( .A1(\seg2/_023_ ), .A2(\seg2/_004_ ), .A3(\seg2/_019_ ), .ZN(\seg2/_035_ ) );
NOR2_X2 \seg2/_086_ ( .A1(\seg2/_034_ ), .A2(\seg2/_035_ ), .ZN(\seg2/_036_ ) );
NAND2_X1 \seg2/_087_ ( .A1(\seg2/_020_ ), .A2(\seg2/_022_ ), .ZN(\seg2/_037_ ) );
NOR2_X4 \seg2/_088_ ( .A1(\seg2/_002_ ), .A2(\seg2/_001_ ), .ZN(\seg2/_038_ ) );
NAND2_X1 \seg2/_089_ ( .A1(\seg2/_026_ ), .A2(\seg2/_038_ ), .ZN(\seg2/_039_ ) );
NAND4_X1 \seg2/_090_ ( .A1(\seg2/_036_ ), .A2(\seg2/_037_ ), .A3(\seg2/_025_ ), .A4(\seg2/_039_ ), .ZN(\seg2/_040_ ) );
NAND2_X1 \seg2/_091_ ( .A1(\seg2/_040_ ), .A2(\seg2/_000_ ), .ZN(\seg2/_007_ ) );
AND2_X1 \seg2/_092_ ( .A1(\seg2/_019_ ), .A2(\seg2/_038_ ), .ZN(\seg2/_041_ ) );
OR4_X4 \seg2/_093_ ( .A1(\seg2/_018_ ), .A2(\seg2/_034_ ), .A3(\seg2/_041_ ), .A4(\seg2/_032_ ), .ZN(\seg2/_042_ ) );
AND2_X1 \seg2/_094_ ( .A1(\seg2/_014_ ), .A2(\seg2/_024_ ), .ZN(\seg2/_043_ ) );
NAND2_X1 \seg2/_095_ ( .A1(\seg2/_043_ ), .A2(\seg2/_031_ ), .ZN(\seg2/_044_ ) );
NAND2_X1 \seg2/_096_ ( .A1(\seg2/_020_ ), .A2(\seg2/_031_ ), .ZN(\seg2/_045_ ) );
NAND3_X1 \seg2/_097_ ( .A1(\seg2/_044_ ), .A2(\seg2/_045_ ), .A3(\seg2/_037_ ), .ZN(\seg2/_046_ ) );
OAI21_X1 \seg2/_098_ ( .A(\seg2/_000_ ), .B1(\seg2/_042_ ), .B2(\seg2/_046_ ), .ZN(\seg2/_008_ ) );
INV_X1 \seg2/_099_ ( .A(\seg2/_043_ ), .ZN(\seg2/_047_ ) );
OAI21_X1 \seg2/_100_ ( .A(\seg2/_044_ ), .B1(\seg2/_047_ ), .B2(\seg2/_033_ ), .ZN(\seg2/_048_ ) );
NAND2_X1 \seg2/_101_ ( .A1(\seg2/_041_ ), .A2(\seg2/_004_ ), .ZN(\seg2/_049_ ) );
NAND2_X1 \seg2/_102_ ( .A1(\seg2/_026_ ), .A2(\seg2/_033_ ), .ZN(\seg2/_050_ ) );
NAND3_X1 \seg2/_103_ ( .A1(\seg2/_023_ ), .A2(\seg2/_004_ ), .A3(\seg2/_014_ ), .ZN(\seg2/_051_ ) );
NAND3_X1 \seg2/_104_ ( .A1(\seg2/_019_ ), .A2(\seg2/_001_ ), .A3(\seg2/_004_ ), .ZN(\seg2/_052_ ) );
NAND4_X1 \seg2/_105_ ( .A1(\seg2/_049_ ), .A2(\seg2/_050_ ), .A3(\seg2/_051_ ), .A4(\seg2/_052_ ), .ZN(\seg2/_053_ ) );
OAI21_X1 \seg2/_106_ ( .A(\seg2/_000_ ), .B1(\seg2/_048_ ), .B2(\seg2/_053_ ), .ZN(\seg2/_009_ ) );
INV_X1 \seg2/_107_ ( .A(\seg2/_021_ ), .ZN(\seg2/_054_ ) );
AOI211_X4 \seg2/_108_ ( .A(\seg2/_005_ ), .B(\seg2/_004_ ), .C1(\seg2/_031_ ), .C2(\seg2/_013_ ), .ZN(\seg2/_055_ ) );
OAI21_X1 \seg2/_109_ ( .A(\seg2/_000_ ), .B1(\seg2/_054_ ), .B2(\seg2/_055_ ), .ZN(\seg2/_010_ ) );
NAND3_X1 \seg2/_110_ ( .A1(\seg2/_014_ ), .A2(\seg2/_030_ ), .A3(\seg2/_024_ ), .ZN(\seg2/_056_ ) );
NOR2_X1 \seg2/_111_ ( .A1(\seg2/_056_ ), .A2(\seg2/_001_ ), .ZN(\seg2/_057_ ) );
OR3_X2 \seg2/_112_ ( .A1(\seg2/_018_ ), .A2(\seg2/_057_ ), .A3(\seg2/_035_ ), .ZN(\seg2/_058_ ) );
AOI211_X4 \seg2/_113_ ( .A(\seg2/_005_ ), .B(\seg2/_004_ ), .C1(\seg2/_023_ ), .C2(\seg2/_003_ ), .ZN(\seg2/_059_ ) );
OAI21_X1 \seg2/_114_ ( .A(\seg2/_000_ ), .B1(\seg2/_058_ ), .B2(\seg2/_059_ ), .ZN(\seg2/_011_ ) );
OAI211_X2 \seg2/_115_ ( .A(\seg2/_036_ ), .B(\seg2/_050_ ), .C1(\seg2/_038_ ), .C2(\seg2/_047_ ), .ZN(\seg2/_060_ ) );
NAND2_X1 \seg2/_116_ ( .A1(\seg2/_060_ ), .A2(\seg2/_000_ ), .ZN(\seg2/_012_ ) );
LOGIC1_X1 \seg2/_117_ ( .Z(\seg2/_061_ ) );
BUF_X1 \seg2/_118_ ( .A(\seg2/_061_ ), .Z(\io_seg_out_2[0] ) );
BUF_X1 \seg2/_119_ ( .A(display_en ), .Z(\seg2/_000_ ) );
BUF_X1 \seg2/_120_ ( .A(_194_ ), .Z(\seg2/_005_ ) );
BUF_X1 \seg2/_121_ ( .A(\seg2_in[1] ), .Z(\seg2/_002_ ) );
BUF_X1 \seg2/_122_ ( .A(\seg2_in[0] ), .Z(\seg2/_001_ ) );
BUF_X1 \seg2/_123_ ( .A(\seg2_in[3] ), .Z(\seg2/_004_ ) );
BUF_X1 \seg2/_124_ ( .A(\seg2_in[2] ), .Z(\seg2/_003_ ) );
BUF_X1 \seg2/_125_ ( .A(\seg2/_006_ ), .Z(\io_seg_out_2[1] ) );
BUF_X1 \seg2/_126_ ( .A(\seg2/_007_ ), .Z(\io_seg_out_2[2] ) );
BUF_X1 \seg2/_127_ ( .A(\seg2/_008_ ), .Z(\io_seg_out_2[3] ) );
BUF_X1 \seg2/_128_ ( .A(\seg2/_009_ ), .Z(\io_seg_out_2[4] ) );
BUF_X1 \seg2/_129_ ( .A(\seg2/_010_ ), .Z(\io_seg_out_2[5] ) );
BUF_X1 \seg2/_130_ ( .A(\seg2/_011_ ), .Z(\io_seg_out_2[6] ) );
BUF_X1 \seg2/_131_ ( .A(\seg2/_012_ ), .Z(\io_seg_out_2[7] ) );
INV_X32 \seg3/_062_ ( .A(\seg3/_003_ ), .ZN(\seg3/_013_ ) );
NOR2_X4 \seg3/_063_ ( .A1(\seg3/_013_ ), .A2(\seg3/_005_ ), .ZN(\seg3/_014_ ) );
AND2_X4 \seg3/_064_ ( .A1(\seg3/_014_ ), .A2(\seg3/_004_ ), .ZN(\seg3/_015_ ) );
INV_X32 \seg3/_065_ ( .A(\seg3/_001_ ), .ZN(\seg3/_016_ ) );
NOR2_X4 \seg3/_066_ ( .A1(\seg3/_016_ ), .A2(\seg3/_002_ ), .ZN(\seg3/_017_ ) );
AND2_X2 \seg3/_067_ ( .A1(\seg3/_015_ ), .A2(\seg3/_017_ ), .ZN(\seg3/_018_ ) );
NOR2_X4 \seg3/_068_ ( .A1(\seg3/_005_ ), .A2(\seg3/_003_ ), .ZN(\seg3/_019_ ) );
AND2_X1 \seg3/_069_ ( .A1(\seg3/_019_ ), .A2(\seg3/_004_ ), .ZN(\seg3/_020_ ) );
NOR2_X2 \seg3/_070_ ( .A1(\seg3/_018_ ), .A2(\seg3/_020_ ), .ZN(\seg3/_021_ ) );
AND2_X4 \seg3/_071_ ( .A1(\seg3/_002_ ), .A2(\seg3/_001_ ), .ZN(\seg3/_022_ ) );
INV_X4 \seg3/_072_ ( .A(\seg3/_022_ ), .ZN(\seg3/_023_ ) );
INV_X32 \seg3/_073_ ( .A(\seg3/_004_ ), .ZN(\seg3/_024_ ) );
NAND3_X1 \seg3/_074_ ( .A1(\seg3/_023_ ), .A2(\seg3/_024_ ), .A3(\seg3/_014_ ), .ZN(\seg3/_025_ ) );
AND2_X4 \seg3/_075_ ( .A1(\seg3/_019_ ), .A2(\seg3/_024_ ), .ZN(\seg3/_026_ ) );
NAND2_X1 \seg3/_076_ ( .A1(\seg3/_026_ ), .A2(\seg3/_022_ ), .ZN(\seg3/_027_ ) );
NAND2_X1 \seg3/_077_ ( .A1(\seg3/_015_ ), .A2(\seg3/_002_ ), .ZN(\seg3/_028_ ) );
NAND4_X1 \seg3/_078_ ( .A1(\seg3/_021_ ), .A2(\seg3/_025_ ), .A3(\seg3/_027_ ), .A4(\seg3/_028_ ), .ZN(\seg3/_029_ ) );
INV_X16 \seg3/_079_ ( .A(\seg3/_002_ ), .ZN(\seg3/_030_ ) );
NOR2_X4 \seg3/_080_ ( .A1(\seg3/_030_ ), .A2(\seg3/_001_ ), .ZN(\seg3/_031_ ) );
AND2_X4 \seg3/_081_ ( .A1(\seg3/_026_ ), .A2(\seg3/_031_ ), .ZN(\seg3/_032_ ) );
OAI21_X1 \seg3/_082_ ( .A(\seg3/_000_ ), .B1(\seg3/_029_ ), .B2(\seg3/_032_ ), .ZN(\seg3/_006_ ) );
INV_X1 \seg3/_083_ ( .A(\seg3/_017_ ), .ZN(\seg3/_033_ ) );
AND2_X4 \seg3/_084_ ( .A1(\seg3/_015_ ), .A2(\seg3/_033_ ), .ZN(\seg3/_034_ ) );
AND3_X2 \seg3/_085_ ( .A1(\seg3/_023_ ), .A2(\seg3/_004_ ), .A3(\seg3/_019_ ), .ZN(\seg3/_035_ ) );
NOR2_X2 \seg3/_086_ ( .A1(\seg3/_034_ ), .A2(\seg3/_035_ ), .ZN(\seg3/_036_ ) );
NAND2_X1 \seg3/_087_ ( .A1(\seg3/_020_ ), .A2(\seg3/_022_ ), .ZN(\seg3/_037_ ) );
NOR2_X4 \seg3/_088_ ( .A1(\seg3/_002_ ), .A2(\seg3/_001_ ), .ZN(\seg3/_038_ ) );
NAND2_X1 \seg3/_089_ ( .A1(\seg3/_026_ ), .A2(\seg3/_038_ ), .ZN(\seg3/_039_ ) );
NAND4_X1 \seg3/_090_ ( .A1(\seg3/_036_ ), .A2(\seg3/_037_ ), .A3(\seg3/_025_ ), .A4(\seg3/_039_ ), .ZN(\seg3/_040_ ) );
NAND2_X1 \seg3/_091_ ( .A1(\seg3/_040_ ), .A2(\seg3/_000_ ), .ZN(\seg3/_007_ ) );
AND2_X1 \seg3/_092_ ( .A1(\seg3/_019_ ), .A2(\seg3/_038_ ), .ZN(\seg3/_041_ ) );
OR4_X4 \seg3/_093_ ( .A1(\seg3/_018_ ), .A2(\seg3/_034_ ), .A3(\seg3/_041_ ), .A4(\seg3/_032_ ), .ZN(\seg3/_042_ ) );
AND2_X1 \seg3/_094_ ( .A1(\seg3/_014_ ), .A2(\seg3/_024_ ), .ZN(\seg3/_043_ ) );
NAND2_X1 \seg3/_095_ ( .A1(\seg3/_043_ ), .A2(\seg3/_031_ ), .ZN(\seg3/_044_ ) );
NAND2_X1 \seg3/_096_ ( .A1(\seg3/_020_ ), .A2(\seg3/_031_ ), .ZN(\seg3/_045_ ) );
NAND3_X1 \seg3/_097_ ( .A1(\seg3/_044_ ), .A2(\seg3/_045_ ), .A3(\seg3/_037_ ), .ZN(\seg3/_046_ ) );
OAI21_X1 \seg3/_098_ ( .A(\seg3/_000_ ), .B1(\seg3/_042_ ), .B2(\seg3/_046_ ), .ZN(\seg3/_008_ ) );
INV_X1 \seg3/_099_ ( .A(\seg3/_043_ ), .ZN(\seg3/_047_ ) );
OAI21_X1 \seg3/_100_ ( .A(\seg3/_044_ ), .B1(\seg3/_047_ ), .B2(\seg3/_033_ ), .ZN(\seg3/_048_ ) );
NAND2_X1 \seg3/_101_ ( .A1(\seg3/_041_ ), .A2(\seg3/_004_ ), .ZN(\seg3/_049_ ) );
NAND2_X1 \seg3/_102_ ( .A1(\seg3/_026_ ), .A2(\seg3/_033_ ), .ZN(\seg3/_050_ ) );
NAND3_X1 \seg3/_103_ ( .A1(\seg3/_023_ ), .A2(\seg3/_004_ ), .A3(\seg3/_014_ ), .ZN(\seg3/_051_ ) );
NAND3_X1 \seg3/_104_ ( .A1(\seg3/_019_ ), .A2(\seg3/_001_ ), .A3(\seg3/_004_ ), .ZN(\seg3/_052_ ) );
NAND4_X1 \seg3/_105_ ( .A1(\seg3/_049_ ), .A2(\seg3/_050_ ), .A3(\seg3/_051_ ), .A4(\seg3/_052_ ), .ZN(\seg3/_053_ ) );
OAI21_X1 \seg3/_106_ ( .A(\seg3/_000_ ), .B1(\seg3/_048_ ), .B2(\seg3/_053_ ), .ZN(\seg3/_009_ ) );
INV_X1 \seg3/_107_ ( .A(\seg3/_021_ ), .ZN(\seg3/_054_ ) );
AOI211_X4 \seg3/_108_ ( .A(\seg3/_005_ ), .B(\seg3/_004_ ), .C1(\seg3/_031_ ), .C2(\seg3/_013_ ), .ZN(\seg3/_055_ ) );
OAI21_X1 \seg3/_109_ ( .A(\seg3/_000_ ), .B1(\seg3/_054_ ), .B2(\seg3/_055_ ), .ZN(\seg3/_010_ ) );
NAND3_X1 \seg3/_110_ ( .A1(\seg3/_014_ ), .A2(\seg3/_030_ ), .A3(\seg3/_024_ ), .ZN(\seg3/_056_ ) );
NOR2_X1 \seg3/_111_ ( .A1(\seg3/_056_ ), .A2(\seg3/_001_ ), .ZN(\seg3/_057_ ) );
OR3_X2 \seg3/_112_ ( .A1(\seg3/_018_ ), .A2(\seg3/_057_ ), .A3(\seg3/_035_ ), .ZN(\seg3/_058_ ) );
AOI211_X4 \seg3/_113_ ( .A(\seg3/_005_ ), .B(\seg3/_004_ ), .C1(\seg3/_023_ ), .C2(\seg3/_003_ ), .ZN(\seg3/_059_ ) );
OAI21_X1 \seg3/_114_ ( .A(\seg3/_000_ ), .B1(\seg3/_058_ ), .B2(\seg3/_059_ ), .ZN(\seg3/_011_ ) );
OAI211_X2 \seg3/_115_ ( .A(\seg3/_036_ ), .B(\seg3/_050_ ), .C1(\seg3/_038_ ), .C2(\seg3/_047_ ), .ZN(\seg3/_060_ ) );
NAND2_X1 \seg3/_116_ ( .A1(\seg3/_060_ ), .A2(\seg3/_000_ ), .ZN(\seg3/_012_ ) );
LOGIC1_X1 \seg3/_117_ ( .Z(\seg3/_061_ ) );
BUF_X1 \seg3/_118_ ( .A(\seg3/_061_ ), .Z(\io_seg_out_3[0] ) );
BUF_X1 \seg3/_119_ ( .A(display_en ), .Z(\seg3/_000_ ) );
BUF_X1 \seg3/_120_ ( .A(_194_ ), .Z(\seg3/_005_ ) );
BUF_X1 \seg3/_121_ ( .A(\seg3_in[1] ), .Z(\seg3/_002_ ) );
BUF_X1 \seg3/_122_ ( .A(\seg3_in[0] ), .Z(\seg3/_001_ ) );
BUF_X1 \seg3/_123_ ( .A(\seg3_in[3] ), .Z(\seg3/_004_ ) );
BUF_X1 \seg3/_124_ ( .A(\seg3_in[2] ), .Z(\seg3/_003_ ) );
BUF_X1 \seg3/_125_ ( .A(\seg3/_006_ ), .Z(\io_seg_out_3[1] ) );
BUF_X1 \seg3/_126_ ( .A(\seg3/_007_ ), .Z(\io_seg_out_3[2] ) );
BUF_X1 \seg3/_127_ ( .A(\seg3/_008_ ), .Z(\io_seg_out_3[3] ) );
BUF_X1 \seg3/_128_ ( .A(\seg3/_009_ ), .Z(\io_seg_out_3[4] ) );
BUF_X1 \seg3/_129_ ( .A(\seg3/_010_ ), .Z(\io_seg_out_3[5] ) );
BUF_X1 \seg3/_130_ ( .A(\seg3/_011_ ), .Z(\io_seg_out_3[6] ) );
BUF_X1 \seg3/_131_ ( .A(\seg3/_012_ ), .Z(\io_seg_out_3[7] ) );
INV_X32 \seg4/_062_ ( .A(\seg4/_003_ ), .ZN(\seg4/_013_ ) );
NOR2_X4 \seg4/_063_ ( .A1(\seg4/_013_ ), .A2(\seg4/_005_ ), .ZN(\seg4/_014_ ) );
AND2_X4 \seg4/_064_ ( .A1(\seg4/_014_ ), .A2(\seg4/_004_ ), .ZN(\seg4/_015_ ) );
INV_X32 \seg4/_065_ ( .A(\seg4/_001_ ), .ZN(\seg4/_016_ ) );
NOR2_X4 \seg4/_066_ ( .A1(\seg4/_016_ ), .A2(\seg4/_002_ ), .ZN(\seg4/_017_ ) );
AND2_X2 \seg4/_067_ ( .A1(\seg4/_015_ ), .A2(\seg4/_017_ ), .ZN(\seg4/_018_ ) );
NOR2_X4 \seg4/_068_ ( .A1(\seg4/_005_ ), .A2(\seg4/_003_ ), .ZN(\seg4/_019_ ) );
AND2_X1 \seg4/_069_ ( .A1(\seg4/_019_ ), .A2(\seg4/_004_ ), .ZN(\seg4/_020_ ) );
NOR2_X2 \seg4/_070_ ( .A1(\seg4/_018_ ), .A2(\seg4/_020_ ), .ZN(\seg4/_021_ ) );
AND2_X4 \seg4/_071_ ( .A1(\seg4/_002_ ), .A2(\seg4/_001_ ), .ZN(\seg4/_022_ ) );
INV_X4 \seg4/_072_ ( .A(\seg4/_022_ ), .ZN(\seg4/_023_ ) );
INV_X32 \seg4/_073_ ( .A(\seg4/_004_ ), .ZN(\seg4/_024_ ) );
NAND3_X1 \seg4/_074_ ( .A1(\seg4/_023_ ), .A2(\seg4/_024_ ), .A3(\seg4/_014_ ), .ZN(\seg4/_025_ ) );
AND2_X4 \seg4/_075_ ( .A1(\seg4/_019_ ), .A2(\seg4/_024_ ), .ZN(\seg4/_026_ ) );
NAND2_X1 \seg4/_076_ ( .A1(\seg4/_026_ ), .A2(\seg4/_022_ ), .ZN(\seg4/_027_ ) );
NAND2_X1 \seg4/_077_ ( .A1(\seg4/_015_ ), .A2(\seg4/_002_ ), .ZN(\seg4/_028_ ) );
NAND4_X1 \seg4/_078_ ( .A1(\seg4/_021_ ), .A2(\seg4/_025_ ), .A3(\seg4/_027_ ), .A4(\seg4/_028_ ), .ZN(\seg4/_029_ ) );
INV_X16 \seg4/_079_ ( .A(\seg4/_002_ ), .ZN(\seg4/_030_ ) );
NOR2_X4 \seg4/_080_ ( .A1(\seg4/_030_ ), .A2(\seg4/_001_ ), .ZN(\seg4/_031_ ) );
AND2_X4 \seg4/_081_ ( .A1(\seg4/_026_ ), .A2(\seg4/_031_ ), .ZN(\seg4/_032_ ) );
OAI21_X1 \seg4/_082_ ( .A(\seg4/_000_ ), .B1(\seg4/_029_ ), .B2(\seg4/_032_ ), .ZN(\seg4/_006_ ) );
INV_X1 \seg4/_083_ ( .A(\seg4/_017_ ), .ZN(\seg4/_033_ ) );
AND2_X4 \seg4/_084_ ( .A1(\seg4/_015_ ), .A2(\seg4/_033_ ), .ZN(\seg4/_034_ ) );
AND3_X2 \seg4/_085_ ( .A1(\seg4/_023_ ), .A2(\seg4/_004_ ), .A3(\seg4/_019_ ), .ZN(\seg4/_035_ ) );
NOR2_X2 \seg4/_086_ ( .A1(\seg4/_034_ ), .A2(\seg4/_035_ ), .ZN(\seg4/_036_ ) );
NAND2_X1 \seg4/_087_ ( .A1(\seg4/_020_ ), .A2(\seg4/_022_ ), .ZN(\seg4/_037_ ) );
NOR2_X4 \seg4/_088_ ( .A1(\seg4/_002_ ), .A2(\seg4/_001_ ), .ZN(\seg4/_038_ ) );
NAND2_X1 \seg4/_089_ ( .A1(\seg4/_026_ ), .A2(\seg4/_038_ ), .ZN(\seg4/_039_ ) );
NAND4_X1 \seg4/_090_ ( .A1(\seg4/_036_ ), .A2(\seg4/_037_ ), .A3(\seg4/_025_ ), .A4(\seg4/_039_ ), .ZN(\seg4/_040_ ) );
NAND2_X1 \seg4/_091_ ( .A1(\seg4/_040_ ), .A2(\seg4/_000_ ), .ZN(\seg4/_007_ ) );
AND2_X1 \seg4/_092_ ( .A1(\seg4/_019_ ), .A2(\seg4/_038_ ), .ZN(\seg4/_041_ ) );
OR4_X4 \seg4/_093_ ( .A1(\seg4/_018_ ), .A2(\seg4/_034_ ), .A3(\seg4/_041_ ), .A4(\seg4/_032_ ), .ZN(\seg4/_042_ ) );
AND2_X1 \seg4/_094_ ( .A1(\seg4/_014_ ), .A2(\seg4/_024_ ), .ZN(\seg4/_043_ ) );
NAND2_X1 \seg4/_095_ ( .A1(\seg4/_043_ ), .A2(\seg4/_031_ ), .ZN(\seg4/_044_ ) );
NAND2_X1 \seg4/_096_ ( .A1(\seg4/_020_ ), .A2(\seg4/_031_ ), .ZN(\seg4/_045_ ) );
NAND3_X1 \seg4/_097_ ( .A1(\seg4/_044_ ), .A2(\seg4/_045_ ), .A3(\seg4/_037_ ), .ZN(\seg4/_046_ ) );
OAI21_X1 \seg4/_098_ ( .A(\seg4/_000_ ), .B1(\seg4/_042_ ), .B2(\seg4/_046_ ), .ZN(\seg4/_008_ ) );
INV_X1 \seg4/_099_ ( .A(\seg4/_043_ ), .ZN(\seg4/_047_ ) );
OAI21_X1 \seg4/_100_ ( .A(\seg4/_044_ ), .B1(\seg4/_047_ ), .B2(\seg4/_033_ ), .ZN(\seg4/_048_ ) );
NAND2_X1 \seg4/_101_ ( .A1(\seg4/_041_ ), .A2(\seg4/_004_ ), .ZN(\seg4/_049_ ) );
NAND2_X1 \seg4/_102_ ( .A1(\seg4/_026_ ), .A2(\seg4/_033_ ), .ZN(\seg4/_050_ ) );
NAND3_X1 \seg4/_103_ ( .A1(\seg4/_023_ ), .A2(\seg4/_004_ ), .A3(\seg4/_014_ ), .ZN(\seg4/_051_ ) );
NAND3_X1 \seg4/_104_ ( .A1(\seg4/_019_ ), .A2(\seg4/_001_ ), .A3(\seg4/_004_ ), .ZN(\seg4/_052_ ) );
NAND4_X1 \seg4/_105_ ( .A1(\seg4/_049_ ), .A2(\seg4/_050_ ), .A3(\seg4/_051_ ), .A4(\seg4/_052_ ), .ZN(\seg4/_053_ ) );
OAI21_X1 \seg4/_106_ ( .A(\seg4/_000_ ), .B1(\seg4/_048_ ), .B2(\seg4/_053_ ), .ZN(\seg4/_009_ ) );
INV_X1 \seg4/_107_ ( .A(\seg4/_021_ ), .ZN(\seg4/_054_ ) );
AOI211_X4 \seg4/_108_ ( .A(\seg4/_005_ ), .B(\seg4/_004_ ), .C1(\seg4/_031_ ), .C2(\seg4/_013_ ), .ZN(\seg4/_055_ ) );
OAI21_X1 \seg4/_109_ ( .A(\seg4/_000_ ), .B1(\seg4/_054_ ), .B2(\seg4/_055_ ), .ZN(\seg4/_010_ ) );
NAND3_X1 \seg4/_110_ ( .A1(\seg4/_014_ ), .A2(\seg4/_030_ ), .A3(\seg4/_024_ ), .ZN(\seg4/_056_ ) );
NOR2_X1 \seg4/_111_ ( .A1(\seg4/_056_ ), .A2(\seg4/_001_ ), .ZN(\seg4/_057_ ) );
OR3_X2 \seg4/_112_ ( .A1(\seg4/_018_ ), .A2(\seg4/_057_ ), .A3(\seg4/_035_ ), .ZN(\seg4/_058_ ) );
AOI211_X4 \seg4/_113_ ( .A(\seg4/_005_ ), .B(\seg4/_004_ ), .C1(\seg4/_023_ ), .C2(\seg4/_003_ ), .ZN(\seg4/_059_ ) );
OAI21_X1 \seg4/_114_ ( .A(\seg4/_000_ ), .B1(\seg4/_058_ ), .B2(\seg4/_059_ ), .ZN(\seg4/_011_ ) );
OAI211_X2 \seg4/_115_ ( .A(\seg4/_036_ ), .B(\seg4/_050_ ), .C1(\seg4/_038_ ), .C2(\seg4/_047_ ), .ZN(\seg4/_060_ ) );
NAND2_X1 \seg4/_116_ ( .A1(\seg4/_060_ ), .A2(\seg4/_000_ ), .ZN(\seg4/_012_ ) );
LOGIC1_X1 \seg4/_117_ ( .Z(\seg4/_061_ ) );
BUF_X1 \seg4/_118_ ( .A(\seg4/_061_ ), .Z(\io_seg_out_4[0] ) );
BUF_X1 \seg4/_119_ ( .A(_193_ ), .Z(\seg4/_000_ ) );
BUF_X1 \seg4/_120_ ( .A(_194_ ), .Z(\seg4/_005_ ) );
BUF_X1 \seg4/_121_ ( .A(\counter_io_ones[1] ), .Z(\seg4/_002_ ) );
BUF_X1 \seg4/_122_ ( .A(\counter_io_ones[0] ), .Z(\seg4/_001_ ) );
BUF_X1 \seg4/_123_ ( .A(\counter_io_ones[3] ), .Z(\seg4/_004_ ) );
BUF_X1 \seg4/_124_ ( .A(\counter_io_ones[2] ), .Z(\seg4/_003_ ) );
BUF_X1 \seg4/_125_ ( .A(\seg4/_006_ ), .Z(\io_seg_out_4[1] ) );
BUF_X1 \seg4/_126_ ( .A(\seg4/_007_ ), .Z(\io_seg_out_4[2] ) );
BUF_X1 \seg4/_127_ ( .A(\seg4/_008_ ), .Z(\io_seg_out_4[3] ) );
BUF_X1 \seg4/_128_ ( .A(\seg4/_009_ ), .Z(\io_seg_out_4[4] ) );
BUF_X1 \seg4/_129_ ( .A(\seg4/_010_ ), .Z(\io_seg_out_4[5] ) );
BUF_X1 \seg4/_130_ ( .A(\seg4/_011_ ), .Z(\io_seg_out_4[6] ) );
BUF_X1 \seg4/_131_ ( .A(\seg4/_012_ ), .Z(\io_seg_out_4[7] ) );
INV_X32 \seg5/_062_ ( .A(\seg5/_003_ ), .ZN(\seg5/_013_ ) );
NOR2_X4 \seg5/_063_ ( .A1(\seg5/_013_ ), .A2(\seg5/_005_ ), .ZN(\seg5/_014_ ) );
AND2_X4 \seg5/_064_ ( .A1(\seg5/_014_ ), .A2(\seg5/_004_ ), .ZN(\seg5/_015_ ) );
INV_X32 \seg5/_065_ ( .A(\seg5/_001_ ), .ZN(\seg5/_016_ ) );
NOR2_X4 \seg5/_066_ ( .A1(\seg5/_016_ ), .A2(\seg5/_002_ ), .ZN(\seg5/_017_ ) );
AND2_X2 \seg5/_067_ ( .A1(\seg5/_015_ ), .A2(\seg5/_017_ ), .ZN(\seg5/_018_ ) );
NOR2_X4 \seg5/_068_ ( .A1(\seg5/_005_ ), .A2(\seg5/_003_ ), .ZN(\seg5/_019_ ) );
AND2_X1 \seg5/_069_ ( .A1(\seg5/_019_ ), .A2(\seg5/_004_ ), .ZN(\seg5/_020_ ) );
NOR2_X2 \seg5/_070_ ( .A1(\seg5/_018_ ), .A2(\seg5/_020_ ), .ZN(\seg5/_021_ ) );
AND2_X4 \seg5/_071_ ( .A1(\seg5/_002_ ), .A2(\seg5/_001_ ), .ZN(\seg5/_022_ ) );
INV_X4 \seg5/_072_ ( .A(\seg5/_022_ ), .ZN(\seg5/_023_ ) );
INV_X32 \seg5/_073_ ( .A(\seg5/_004_ ), .ZN(\seg5/_024_ ) );
NAND3_X1 \seg5/_074_ ( .A1(\seg5/_023_ ), .A2(\seg5/_024_ ), .A3(\seg5/_014_ ), .ZN(\seg5/_025_ ) );
AND2_X4 \seg5/_075_ ( .A1(\seg5/_019_ ), .A2(\seg5/_024_ ), .ZN(\seg5/_026_ ) );
NAND2_X1 \seg5/_076_ ( .A1(\seg5/_026_ ), .A2(\seg5/_022_ ), .ZN(\seg5/_027_ ) );
NAND2_X1 \seg5/_077_ ( .A1(\seg5/_015_ ), .A2(\seg5/_002_ ), .ZN(\seg5/_028_ ) );
NAND4_X1 \seg5/_078_ ( .A1(\seg5/_021_ ), .A2(\seg5/_025_ ), .A3(\seg5/_027_ ), .A4(\seg5/_028_ ), .ZN(\seg5/_029_ ) );
INV_X16 \seg5/_079_ ( .A(\seg5/_002_ ), .ZN(\seg5/_030_ ) );
NOR2_X4 \seg5/_080_ ( .A1(\seg5/_030_ ), .A2(\seg5/_001_ ), .ZN(\seg5/_031_ ) );
AND2_X4 \seg5/_081_ ( .A1(\seg5/_026_ ), .A2(\seg5/_031_ ), .ZN(\seg5/_032_ ) );
OAI21_X1 \seg5/_082_ ( .A(\seg5/_000_ ), .B1(\seg5/_029_ ), .B2(\seg5/_032_ ), .ZN(\seg5/_006_ ) );
INV_X1 \seg5/_083_ ( .A(\seg5/_017_ ), .ZN(\seg5/_033_ ) );
AND2_X4 \seg5/_084_ ( .A1(\seg5/_015_ ), .A2(\seg5/_033_ ), .ZN(\seg5/_034_ ) );
AND3_X2 \seg5/_085_ ( .A1(\seg5/_023_ ), .A2(\seg5/_004_ ), .A3(\seg5/_019_ ), .ZN(\seg5/_035_ ) );
NOR2_X2 \seg5/_086_ ( .A1(\seg5/_034_ ), .A2(\seg5/_035_ ), .ZN(\seg5/_036_ ) );
NAND2_X1 \seg5/_087_ ( .A1(\seg5/_020_ ), .A2(\seg5/_022_ ), .ZN(\seg5/_037_ ) );
NOR2_X4 \seg5/_088_ ( .A1(\seg5/_002_ ), .A2(\seg5/_001_ ), .ZN(\seg5/_038_ ) );
NAND2_X1 \seg5/_089_ ( .A1(\seg5/_026_ ), .A2(\seg5/_038_ ), .ZN(\seg5/_039_ ) );
NAND4_X1 \seg5/_090_ ( .A1(\seg5/_036_ ), .A2(\seg5/_037_ ), .A3(\seg5/_025_ ), .A4(\seg5/_039_ ), .ZN(\seg5/_040_ ) );
NAND2_X1 \seg5/_091_ ( .A1(\seg5/_040_ ), .A2(\seg5/_000_ ), .ZN(\seg5/_007_ ) );
AND2_X1 \seg5/_092_ ( .A1(\seg5/_019_ ), .A2(\seg5/_038_ ), .ZN(\seg5/_041_ ) );
OR4_X4 \seg5/_093_ ( .A1(\seg5/_018_ ), .A2(\seg5/_034_ ), .A3(\seg5/_041_ ), .A4(\seg5/_032_ ), .ZN(\seg5/_042_ ) );
AND2_X1 \seg5/_094_ ( .A1(\seg5/_014_ ), .A2(\seg5/_024_ ), .ZN(\seg5/_043_ ) );
NAND2_X1 \seg5/_095_ ( .A1(\seg5/_043_ ), .A2(\seg5/_031_ ), .ZN(\seg5/_044_ ) );
NAND2_X1 \seg5/_096_ ( .A1(\seg5/_020_ ), .A2(\seg5/_031_ ), .ZN(\seg5/_045_ ) );
NAND3_X1 \seg5/_097_ ( .A1(\seg5/_044_ ), .A2(\seg5/_045_ ), .A3(\seg5/_037_ ), .ZN(\seg5/_046_ ) );
OAI21_X1 \seg5/_098_ ( .A(\seg5/_000_ ), .B1(\seg5/_042_ ), .B2(\seg5/_046_ ), .ZN(\seg5/_008_ ) );
INV_X1 \seg5/_099_ ( .A(\seg5/_043_ ), .ZN(\seg5/_047_ ) );
OAI21_X1 \seg5/_100_ ( .A(\seg5/_044_ ), .B1(\seg5/_047_ ), .B2(\seg5/_033_ ), .ZN(\seg5/_048_ ) );
NAND2_X1 \seg5/_101_ ( .A1(\seg5/_041_ ), .A2(\seg5/_004_ ), .ZN(\seg5/_049_ ) );
NAND2_X1 \seg5/_102_ ( .A1(\seg5/_026_ ), .A2(\seg5/_033_ ), .ZN(\seg5/_050_ ) );
NAND3_X1 \seg5/_103_ ( .A1(\seg5/_023_ ), .A2(\seg5/_004_ ), .A3(\seg5/_014_ ), .ZN(\seg5/_051_ ) );
NAND3_X1 \seg5/_104_ ( .A1(\seg5/_019_ ), .A2(\seg5/_001_ ), .A3(\seg5/_004_ ), .ZN(\seg5/_052_ ) );
NAND4_X1 \seg5/_105_ ( .A1(\seg5/_049_ ), .A2(\seg5/_050_ ), .A3(\seg5/_051_ ), .A4(\seg5/_052_ ), .ZN(\seg5/_053_ ) );
OAI21_X1 \seg5/_106_ ( .A(\seg5/_000_ ), .B1(\seg5/_048_ ), .B2(\seg5/_053_ ), .ZN(\seg5/_009_ ) );
INV_X1 \seg5/_107_ ( .A(\seg5/_021_ ), .ZN(\seg5/_054_ ) );
AOI211_X4 \seg5/_108_ ( .A(\seg5/_005_ ), .B(\seg5/_004_ ), .C1(\seg5/_031_ ), .C2(\seg5/_013_ ), .ZN(\seg5/_055_ ) );
OAI21_X1 \seg5/_109_ ( .A(\seg5/_000_ ), .B1(\seg5/_054_ ), .B2(\seg5/_055_ ), .ZN(\seg5/_010_ ) );
NAND3_X1 \seg5/_110_ ( .A1(\seg5/_014_ ), .A2(\seg5/_030_ ), .A3(\seg5/_024_ ), .ZN(\seg5/_056_ ) );
NOR2_X1 \seg5/_111_ ( .A1(\seg5/_056_ ), .A2(\seg5/_001_ ), .ZN(\seg5/_057_ ) );
OR3_X2 \seg5/_112_ ( .A1(\seg5/_018_ ), .A2(\seg5/_057_ ), .A3(\seg5/_035_ ), .ZN(\seg5/_058_ ) );
AOI211_X4 \seg5/_113_ ( .A(\seg5/_005_ ), .B(\seg5/_004_ ), .C1(\seg5/_023_ ), .C2(\seg5/_003_ ), .ZN(\seg5/_059_ ) );
OAI21_X1 \seg5/_114_ ( .A(\seg5/_000_ ), .B1(\seg5/_058_ ), .B2(\seg5/_059_ ), .ZN(\seg5/_011_ ) );
OAI211_X2 \seg5/_115_ ( .A(\seg5/_036_ ), .B(\seg5/_050_ ), .C1(\seg5/_038_ ), .C2(\seg5/_047_ ), .ZN(\seg5/_060_ ) );
NAND2_X1 \seg5/_116_ ( .A1(\seg5/_060_ ), .A2(\seg5/_000_ ), .ZN(\seg5/_012_ ) );
LOGIC1_X1 \seg5/_117_ ( .Z(\seg5/_061_ ) );
BUF_X1 \seg5/_118_ ( .A(\seg5/_061_ ), .Z(\io_seg_out_5[0] ) );
BUF_X1 \seg5/_119_ ( .A(_193_ ), .Z(\seg5/_000_ ) );
BUF_X1 \seg5/_120_ ( .A(_194_ ), .Z(\seg5/_005_ ) );
BUF_X1 \seg5/_121_ ( .A(\counter_io_tens[1] ), .Z(\seg5/_002_ ) );
BUF_X1 \seg5/_122_ ( .A(\counter_io_tens[0] ), .Z(\seg5/_001_ ) );
BUF_X1 \seg5/_123_ ( .A(\counter_io_tens[3] ), .Z(\seg5/_004_ ) );
BUF_X1 \seg5/_124_ ( .A(\counter_io_tens[2] ), .Z(\seg5/_003_ ) );
BUF_X1 \seg5/_125_ ( .A(\seg5/_006_ ), .Z(\io_seg_out_5[1] ) );
BUF_X1 \seg5/_126_ ( .A(\seg5/_007_ ), .Z(\io_seg_out_5[2] ) );
BUF_X1 \seg5/_127_ ( .A(\seg5/_008_ ), .Z(\io_seg_out_5[3] ) );
BUF_X1 \seg5/_128_ ( .A(\seg5/_009_ ), .Z(\io_seg_out_5[4] ) );
BUF_X1 \seg5/_129_ ( .A(\seg5/_010_ ), .Z(\io_seg_out_5[5] ) );
BUF_X1 \seg5/_130_ ( .A(\seg5/_011_ ), .Z(\io_seg_out_5[6] ) );
BUF_X1 \seg5/_131_ ( .A(\seg5/_012_ ), .Z(\io_seg_out_5[7] ) );

endmodule
