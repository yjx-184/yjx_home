//Generate the verilog at 2025-02-27T14:39:44
module ps2_top (
clk,
clrn,
overflow,
ps2_clk,
ps2_data,
seg_out_0,
seg_out_1,
seg_out_2,
seg_out_3,
seg_out_4,
seg_out_5
);

input clk ;
input clrn ;
output overflow ;
input ps2_clk ;
input ps2_data ;
output [7:0] seg_out_0 ;
output [7:0] seg_out_1 ;
output [7:0] seg_out_2 ;
output [7:0] seg_out_3 ;
output [7:0] seg_out_4 ;
output [7:0] seg_out_5 ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire en ;
wire key_release ;
wire nextdata_n ;
wire ready ;
wire ready_d1 ;
wire \u0_ps2_kb/_0000_ ;
wire \u0_ps2_kb/_0001_ ;
wire \u0_ps2_kb/_0002_ ;
wire \u0_ps2_kb/_0003_ ;
wire \u0_ps2_kb/_0004_ ;
wire \u0_ps2_kb/_0005_ ;
wire \u0_ps2_kb/_0006_ ;
wire \u0_ps2_kb/_0007_ ;
wire \u0_ps2_kb/_0008_ ;
wire \u0_ps2_kb/_0009_ ;
wire \u0_ps2_kb/_0010_ ;
wire \u0_ps2_kb/_0011_ ;
wire \u0_ps2_kb/_0012_ ;
wire \u0_ps2_kb/_0013_ ;
wire \u0_ps2_kb/_0014_ ;
wire \u0_ps2_kb/_0015_ ;
wire \u0_ps2_kb/_0016_ ;
wire \u0_ps2_kb/_0017_ ;
wire \u0_ps2_kb/_0018_ ;
wire \u0_ps2_kb/_0019_ ;
wire \u0_ps2_kb/_0020_ ;
wire \u0_ps2_kb/_0021_ ;
wire \u0_ps2_kb/_0022_ ;
wire \u0_ps2_kb/_0023_ ;
wire \u0_ps2_kb/_0024_ ;
wire \u0_ps2_kb/_0025_ ;
wire \u0_ps2_kb/_0026_ ;
wire \u0_ps2_kb/_0027_ ;
wire \u0_ps2_kb/_0028_ ;
wire \u0_ps2_kb/_0029_ ;
wire \u0_ps2_kb/_0030_ ;
wire \u0_ps2_kb/_0031_ ;
wire \u0_ps2_kb/_0032_ ;
wire \u0_ps2_kb/_0033_ ;
wire \u0_ps2_kb/_0034_ ;
wire \u0_ps2_kb/_0035_ ;
wire \u0_ps2_kb/_0036_ ;
wire \u0_ps2_kb/_0037_ ;
wire \u0_ps2_kb/_0038_ ;
wire \u0_ps2_kb/_0039_ ;
wire \u0_ps2_kb/_0040_ ;
wire \u0_ps2_kb/_0041_ ;
wire \u0_ps2_kb/_0042_ ;
wire \u0_ps2_kb/_0043_ ;
wire \u0_ps2_kb/_0044_ ;
wire \u0_ps2_kb/_0045_ ;
wire \u0_ps2_kb/_0046_ ;
wire \u0_ps2_kb/_0047_ ;
wire \u0_ps2_kb/_0048_ ;
wire \u0_ps2_kb/_0049_ ;
wire \u0_ps2_kb/_0050_ ;
wire \u0_ps2_kb/_0051_ ;
wire \u0_ps2_kb/_0052_ ;
wire \u0_ps2_kb/_0053_ ;
wire \u0_ps2_kb/_0054_ ;
wire \u0_ps2_kb/_0055_ ;
wire \u0_ps2_kb/_0056_ ;
wire \u0_ps2_kb/_0057_ ;
wire \u0_ps2_kb/_0058_ ;
wire \u0_ps2_kb/_0059_ ;
wire \u0_ps2_kb/_0060_ ;
wire \u0_ps2_kb/_0061_ ;
wire \u0_ps2_kb/_0062_ ;
wire \u0_ps2_kb/_0063_ ;
wire \u0_ps2_kb/_0064_ ;
wire \u0_ps2_kb/_0065_ ;
wire \u0_ps2_kb/_0066_ ;
wire \u0_ps2_kb/_0067_ ;
wire \u0_ps2_kb/_0068_ ;
wire \u0_ps2_kb/_0069_ ;
wire \u0_ps2_kb/_0070_ ;
wire \u0_ps2_kb/_0071_ ;
wire \u0_ps2_kb/_0072_ ;
wire \u0_ps2_kb/_0073_ ;
wire \u0_ps2_kb/_0074_ ;
wire \u0_ps2_kb/_0075_ ;
wire \u0_ps2_kb/_0076_ ;
wire \u0_ps2_kb/_0077_ ;
wire \u0_ps2_kb/_0078_ ;
wire \u0_ps2_kb/_0079_ ;
wire \u0_ps2_kb/_0080_ ;
wire \u0_ps2_kb/_0081_ ;
wire \u0_ps2_kb/_0082_ ;
wire \u0_ps2_kb/_0083_ ;
wire \u0_ps2_kb/_0084_ ;
wire \u0_ps2_kb/_0085_ ;
wire \u0_ps2_kb/_0086_ ;
wire \u0_ps2_kb/_0087_ ;
wire \u0_ps2_kb/_0088_ ;
wire \u0_ps2_kb/_0089_ ;
wire \u0_ps2_kb/_0090_ ;
wire \u0_ps2_kb/_0091_ ;
wire \u0_ps2_kb/_0092_ ;
wire \u0_ps2_kb/_0093_ ;
wire \u0_ps2_kb/_0094_ ;
wire \u0_ps2_kb/_0095_ ;
wire \u0_ps2_kb/_0096_ ;
wire \u0_ps2_kb/_0097_ ;
wire \u0_ps2_kb/_0098_ ;
wire \u0_ps2_kb/_0099_ ;
wire \u0_ps2_kb/_0100_ ;
wire \u0_ps2_kb/_0101_ ;
wire \u0_ps2_kb/_0102_ ;
wire \u0_ps2_kb/_0103_ ;
wire \u0_ps2_kb/_0104_ ;
wire \u0_ps2_kb/_0105_ ;
wire \u0_ps2_kb/_0106_ ;
wire \u0_ps2_kb/_0107_ ;
wire \u0_ps2_kb/_0108_ ;
wire \u0_ps2_kb/_0109_ ;
wire \u0_ps2_kb/_0110_ ;
wire \u0_ps2_kb/_0111_ ;
wire \u0_ps2_kb/_0112_ ;
wire \u0_ps2_kb/_0113_ ;
wire \u0_ps2_kb/_0114_ ;
wire \u0_ps2_kb/_0115_ ;
wire \u0_ps2_kb/_0116_ ;
wire \u0_ps2_kb/_0117_ ;
wire \u0_ps2_kb/_0118_ ;
wire \u0_ps2_kb/_0119_ ;
wire \u0_ps2_kb/_0120_ ;
wire \u0_ps2_kb/_0121_ ;
wire \u0_ps2_kb/_0122_ ;
wire \u0_ps2_kb/_0123_ ;
wire \u0_ps2_kb/_0124_ ;
wire \u0_ps2_kb/_0125_ ;
wire \u0_ps2_kb/_0126_ ;
wire \u0_ps2_kb/_0127_ ;
wire \u0_ps2_kb/_0128_ ;
wire \u0_ps2_kb/_0129_ ;
wire \u0_ps2_kb/_0130_ ;
wire \u0_ps2_kb/_0131_ ;
wire \u0_ps2_kb/_0132_ ;
wire \u0_ps2_kb/_0133_ ;
wire \u0_ps2_kb/_0134_ ;
wire \u0_ps2_kb/_0135_ ;
wire \u0_ps2_kb/_0136_ ;
wire \u0_ps2_kb/_0137_ ;
wire \u0_ps2_kb/_0138_ ;
wire \u0_ps2_kb/_0139_ ;
wire \u0_ps2_kb/_0140_ ;
wire \u0_ps2_kb/_0141_ ;
wire \u0_ps2_kb/_0142_ ;
wire \u0_ps2_kb/_0143_ ;
wire \u0_ps2_kb/_0144_ ;
wire \u0_ps2_kb/_0145_ ;
wire \u0_ps2_kb/_0146_ ;
wire \u0_ps2_kb/_0147_ ;
wire \u0_ps2_kb/_0148_ ;
wire \u0_ps2_kb/_0149_ ;
wire \u0_ps2_kb/_0150_ ;
wire \u0_ps2_kb/_0151_ ;
wire \u0_ps2_kb/_0152_ ;
wire \u0_ps2_kb/_0153_ ;
wire \u0_ps2_kb/_0154_ ;
wire \u0_ps2_kb/_0155_ ;
wire \u0_ps2_kb/_0156_ ;
wire \u0_ps2_kb/_0157_ ;
wire \u0_ps2_kb/_0158_ ;
wire \u0_ps2_kb/_0159_ ;
wire \u0_ps2_kb/_0160_ ;
wire \u0_ps2_kb/_0161_ ;
wire \u0_ps2_kb/_0162_ ;
wire \u0_ps2_kb/_0163_ ;
wire \u0_ps2_kb/_0164_ ;
wire \u0_ps2_kb/_0165_ ;
wire \u0_ps2_kb/_0166_ ;
wire \u0_ps2_kb/_0167_ ;
wire \u0_ps2_kb/_0168_ ;
wire \u0_ps2_kb/_0169_ ;
wire \u0_ps2_kb/_0170_ ;
wire \u0_ps2_kb/_0171_ ;
wire \u0_ps2_kb/_0172_ ;
wire \u0_ps2_kb/_0173_ ;
wire \u0_ps2_kb/_0174_ ;
wire \u0_ps2_kb/_0175_ ;
wire \u0_ps2_kb/_0176_ ;
wire \u0_ps2_kb/_0177_ ;
wire \u0_ps2_kb/_0178_ ;
wire \u0_ps2_kb/_0179_ ;
wire \u0_ps2_kb/_0180_ ;
wire \u0_ps2_kb/_0181_ ;
wire \u0_ps2_kb/_0182_ ;
wire \u0_ps2_kb/_0183_ ;
wire \u0_ps2_kb/_0184_ ;
wire \u0_ps2_kb/_0185_ ;
wire \u0_ps2_kb/_0186_ ;
wire \u0_ps2_kb/_0187_ ;
wire \u0_ps2_kb/_0188_ ;
wire \u0_ps2_kb/_0189_ ;
wire \u0_ps2_kb/_0190_ ;
wire \u0_ps2_kb/_0191_ ;
wire \u0_ps2_kb/_0192_ ;
wire \u0_ps2_kb/_0193_ ;
wire \u0_ps2_kb/_0194_ ;
wire \u0_ps2_kb/_0195_ ;
wire \u0_ps2_kb/_0196_ ;
wire \u0_ps2_kb/_0197_ ;
wire \u0_ps2_kb/_0198_ ;
wire \u0_ps2_kb/_0199_ ;
wire \u0_ps2_kb/_0200_ ;
wire \u0_ps2_kb/_0201_ ;
wire \u0_ps2_kb/_0202_ ;
wire \u0_ps2_kb/_0203_ ;
wire \u0_ps2_kb/_0204_ ;
wire \u0_ps2_kb/_0205_ ;
wire \u0_ps2_kb/_0206_ ;
wire \u0_ps2_kb/_0207_ ;
wire \u0_ps2_kb/_0208_ ;
wire \u0_ps2_kb/_0209_ ;
wire \u0_ps2_kb/_0210_ ;
wire \u0_ps2_kb/_0211_ ;
wire \u0_ps2_kb/_0212_ ;
wire \u0_ps2_kb/_0213_ ;
wire \u0_ps2_kb/_0214_ ;
wire \u0_ps2_kb/_0215_ ;
wire \u0_ps2_kb/_0216_ ;
wire \u0_ps2_kb/_0217_ ;
wire \u0_ps2_kb/_0218_ ;
wire \u0_ps2_kb/_0219_ ;
wire \u0_ps2_kb/_0220_ ;
wire \u0_ps2_kb/_0221_ ;
wire \u0_ps2_kb/_0222_ ;
wire \u0_ps2_kb/_0223_ ;
wire \u0_ps2_kb/_0224_ ;
wire \u0_ps2_kb/_0225_ ;
wire \u0_ps2_kb/_0226_ ;
wire \u0_ps2_kb/_0227_ ;
wire \u0_ps2_kb/_0228_ ;
wire \u0_ps2_kb/_0229_ ;
wire \u0_ps2_kb/_0230_ ;
wire \u0_ps2_kb/_0231_ ;
wire \u0_ps2_kb/_0232_ ;
wire \u0_ps2_kb/_0233_ ;
wire \u0_ps2_kb/_0234_ ;
wire \u0_ps2_kb/_0235_ ;
wire \u0_ps2_kb/_0236_ ;
wire \u0_ps2_kb/_0237_ ;
wire \u0_ps2_kb/_0238_ ;
wire \u0_ps2_kb/_0239_ ;
wire \u0_ps2_kb/_0240_ ;
wire \u0_ps2_kb/_0241_ ;
wire \u0_ps2_kb/_0242_ ;
wire \u0_ps2_kb/_0243_ ;
wire \u0_ps2_kb/_0244_ ;
wire \u0_ps2_kb/_0245_ ;
wire \u0_ps2_kb/_0246_ ;
wire \u0_ps2_kb/_0247_ ;
wire \u0_ps2_kb/_0248_ ;
wire \u0_ps2_kb/_0249_ ;
wire \u0_ps2_kb/_0250_ ;
wire \u0_ps2_kb/_0251_ ;
wire \u0_ps2_kb/_0252_ ;
wire \u0_ps2_kb/_0253_ ;
wire \u0_ps2_kb/_0254_ ;
wire \u0_ps2_kb/_0255_ ;
wire \u0_ps2_kb/_0256_ ;
wire \u0_ps2_kb/_0257_ ;
wire \u0_ps2_kb/_0258_ ;
wire \u0_ps2_kb/_0259_ ;
wire \u0_ps2_kb/_0260_ ;
wire \u0_ps2_kb/_0261_ ;
wire \u0_ps2_kb/_0262_ ;
wire \u0_ps2_kb/_0263_ ;
wire \u0_ps2_kb/_0264_ ;
wire \u0_ps2_kb/_0265_ ;
wire \u0_ps2_kb/_0266_ ;
wire \u0_ps2_kb/_0267_ ;
wire \u0_ps2_kb/_0268_ ;
wire \u0_ps2_kb/_0269_ ;
wire \u0_ps2_kb/_0270_ ;
wire \u0_ps2_kb/_0271_ ;
wire \u0_ps2_kb/_0272_ ;
wire \u0_ps2_kb/_0273_ ;
wire \u0_ps2_kb/_0274_ ;
wire \u0_ps2_kb/_0275_ ;
wire \u0_ps2_kb/_0276_ ;
wire \u0_ps2_kb/_0277_ ;
wire \u0_ps2_kb/_0278_ ;
wire \u0_ps2_kb/_0279_ ;
wire \u0_ps2_kb/_0280_ ;
wire \u0_ps2_kb/_0281_ ;
wire \u0_ps2_kb/_0282_ ;
wire \u0_ps2_kb/_0283_ ;
wire \u0_ps2_kb/_0284_ ;
wire \u0_ps2_kb/_0285_ ;
wire \u0_ps2_kb/_0286_ ;
wire \u0_ps2_kb/_0287_ ;
wire \u0_ps2_kb/_0288_ ;
wire \u0_ps2_kb/_0289_ ;
wire \u0_ps2_kb/_0290_ ;
wire \u0_ps2_kb/_0291_ ;
wire \u0_ps2_kb/_0292_ ;
wire \u0_ps2_kb/_0293_ ;
wire \u0_ps2_kb/_0294_ ;
wire \u0_ps2_kb/_0295_ ;
wire \u0_ps2_kb/_0296_ ;
wire \u0_ps2_kb/_0297_ ;
wire \u0_ps2_kb/_0298_ ;
wire \u0_ps2_kb/_0299_ ;
wire \u0_ps2_kb/_0300_ ;
wire \u0_ps2_kb/_0301_ ;
wire \u0_ps2_kb/_0302_ ;
wire \u0_ps2_kb/_0303_ ;
wire \u0_ps2_kb/_0304_ ;
wire \u0_ps2_kb/_0305_ ;
wire \u0_ps2_kb/_0306_ ;
wire \u0_ps2_kb/_0307_ ;
wire \u0_ps2_kb/_0308_ ;
wire \u0_ps2_kb/_0309_ ;
wire \u0_ps2_kb/_0310_ ;
wire \u0_ps2_kb/_0311_ ;
wire \u0_ps2_kb/_0312_ ;
wire \u0_ps2_kb/_0313_ ;
wire \u0_ps2_kb/_0314_ ;
wire \u0_ps2_kb/_0315_ ;
wire \u0_ps2_kb/_0316_ ;
wire \u0_ps2_kb/_0317_ ;
wire \u0_ps2_kb/_0318_ ;
wire \u0_ps2_kb/_0319_ ;
wire \u0_ps2_kb/_0320_ ;
wire \u0_ps2_kb/_0321_ ;
wire \u0_ps2_kb/_0322_ ;
wire \u0_ps2_kb/_0323_ ;
wire \u0_ps2_kb/_0324_ ;
wire \u0_ps2_kb/_0325_ ;
wire \u0_ps2_kb/_0326_ ;
wire \u0_ps2_kb/_0327_ ;
wire \u0_ps2_kb/_0328_ ;
wire \u0_ps2_kb/_0329_ ;
wire \u0_ps2_kb/_0330_ ;
wire \u0_ps2_kb/_0331_ ;
wire \u0_ps2_kb/_0332_ ;
wire \u0_ps2_kb/_0333_ ;
wire \u0_ps2_kb/_0334_ ;
wire \u0_ps2_kb/_0335_ ;
wire \u0_ps2_kb/_0336_ ;
wire \u0_ps2_kb/_0337_ ;
wire \u0_ps2_kb/_0338_ ;
wire \u0_ps2_kb/_0339_ ;
wire \u0_ps2_kb/_0340_ ;
wire \u0_ps2_kb/_0341_ ;
wire \u0_ps2_kb/_0342_ ;
wire \u0_ps2_kb/_0343_ ;
wire \u0_ps2_kb/_0344_ ;
wire \u0_ps2_kb/_0345_ ;
wire \u0_ps2_kb/_0346_ ;
wire \u0_ps2_kb/_0347_ ;
wire \u0_ps2_kb/_0348_ ;
wire \u0_ps2_kb/_0349_ ;
wire \u0_ps2_kb/_0350_ ;
wire \u0_ps2_kb/_0351_ ;
wire \u0_ps2_kb/_0352_ ;
wire \u0_ps2_kb/_0353_ ;
wire \u0_ps2_kb/_0354_ ;
wire \u0_ps2_kb/_0355_ ;
wire \u0_ps2_kb/_0356_ ;
wire \u0_ps2_kb/_0357_ ;
wire \u0_ps2_kb/_0358_ ;
wire \u0_ps2_kb/_0359_ ;
wire \u0_ps2_kb/_0360_ ;
wire \u0_ps2_kb/_0361_ ;
wire \u0_ps2_kb/_0362_ ;
wire \u0_ps2_kb/_0363_ ;
wire \u0_ps2_kb/_0364_ ;
wire \u0_ps2_kb/_0365_ ;
wire \u0_ps2_kb/_0366_ ;
wire \u0_ps2_kb/_0367_ ;
wire \u0_ps2_kb/_0368_ ;
wire \u0_ps2_kb/_0369_ ;
wire \u0_ps2_kb/_0370_ ;
wire \u0_ps2_kb/_0371_ ;
wire \u0_ps2_kb/_0372_ ;
wire \u0_ps2_kb/_0373_ ;
wire \u0_ps2_kb/_0374_ ;
wire \u0_ps2_kb/_0375_ ;
wire \u0_ps2_kb/_0376_ ;
wire \u0_ps2_kb/_0377_ ;
wire \u0_ps2_kb/_0378_ ;
wire \u0_ps2_kb/_0379_ ;
wire \u0_ps2_kb/_0380_ ;
wire \u0_ps2_kb/_0381_ ;
wire \u0_ps2_kb/_0382_ ;
wire \u0_ps2_kb/_0383_ ;
wire \u0_ps2_kb/_0384_ ;
wire \u0_ps2_kb/_0385_ ;
wire \u0_ps2_kb/_0386_ ;
wire \u0_ps2_kb/_0387_ ;
wire \u0_ps2_kb/_0388_ ;
wire \u0_ps2_kb/_0389_ ;
wire \u0_ps2_kb/_0390_ ;
wire \u0_ps2_kb/_0391_ ;
wire \u0_ps2_kb/_0392_ ;
wire \u0_ps2_kb/_0393_ ;
wire \u0_ps2_kb/_0394_ ;
wire \u0_ps2_kb/_0395_ ;
wire \u0_ps2_kb/_0396_ ;
wire \u0_ps2_kb/_0397_ ;
wire \u0_ps2_kb/_0398_ ;
wire \u0_ps2_kb/_0399_ ;
wire \u0_ps2_kb/_0400_ ;
wire \u0_ps2_kb/_0401_ ;
wire \u0_ps2_kb/_0402_ ;
wire \u0_ps2_kb/_0403_ ;
wire \u0_ps2_kb/_0404_ ;
wire \u0_ps2_kb/_0405_ ;
wire \u0_ps2_kb/_0406_ ;
wire \u0_ps2_kb/_0407_ ;
wire \u0_ps2_kb/_0408_ ;
wire \u0_ps2_kb/_0409_ ;
wire \u0_ps2_kb/_0410_ ;
wire \u0_ps2_kb/_0411_ ;
wire \u0_ps2_kb/_0412_ ;
wire \u0_ps2_kb/_0413_ ;
wire \u0_ps2_kb/_0414_ ;
wire \u0_ps2_kb/_0415_ ;
wire \u0_ps2_kb/_0416_ ;
wire \u0_ps2_kb/_0417_ ;
wire \u0_ps2_kb/_0418_ ;
wire \u0_ps2_kb/_0419_ ;
wire \u0_ps2_kb/_0420_ ;
wire \u0_ps2_kb/_0421_ ;
wire \u0_ps2_kb/_0422_ ;
wire \u0_ps2_kb/_0423_ ;
wire \u0_ps2_kb/_0424_ ;
wire \u0_ps2_kb/_0425_ ;
wire \u0_ps2_kb/_0426_ ;
wire \u0_ps2_kb/_0427_ ;
wire \u0_ps2_kb/_0428_ ;
wire \u0_ps2_kb/_0429_ ;
wire \u0_ps2_kb/_0430_ ;
wire \u0_ps2_kb/_0431_ ;
wire \u0_ps2_kb/_0432_ ;
wire \u0_ps2_kb/_0433_ ;
wire \u0_ps2_kb/_0434_ ;
wire \u0_ps2_kb/_0435_ ;
wire \u0_ps2_kb/_0436_ ;
wire \u0_ps2_kb/_0437_ ;
wire \u0_ps2_kb/_0438_ ;
wire \u0_ps2_kb/_0439_ ;
wire \u0_ps2_kb/_0440_ ;
wire \u0_ps2_kb/_0441_ ;
wire \u0_ps2_kb/_0442_ ;
wire \u0_ps2_kb/_0443_ ;
wire \u0_ps2_kb/_0444_ ;
wire \u0_ps2_kb/_0445_ ;
wire \u0_ps2_kb/_0446_ ;
wire \u0_ps2_kb/_0447_ ;
wire \u0_ps2_kb/_0448_ ;
wire \u0_ps2_kb/_0449_ ;
wire \u0_ps2_kb/_0450_ ;
wire \u0_ps2_kb/_0451_ ;
wire \u0_ps2_kb/_0452_ ;
wire \u0_ps2_kb/_0453_ ;
wire \u0_ps2_kb/_0454_ ;
wire \u0_ps2_kb/_0455_ ;
wire \u0_ps2_kb/_0456_ ;
wire \u0_ps2_kb/_0457_ ;
wire \u0_ps2_kb/_0458_ ;
wire \u0_ps2_kb/_0459_ ;
wire \u0_ps2_kb/_0460_ ;
wire \u0_ps2_kb/_0461_ ;
wire \u0_ps2_kb/_0462_ ;
wire \u0_ps2_kb/_0463_ ;
wire \u0_ps2_kb/_0464_ ;
wire \u0_ps2_kb/_0465_ ;
wire \u0_ps2_kb/_0466_ ;
wire \u0_ps2_kb/_0467_ ;
wire \u0_ps2_kb/_0468_ ;
wire \u0_ps2_kb/_0469_ ;
wire \u0_ps2_kb/_0470_ ;
wire \u0_ps2_kb/_0471_ ;
wire \u0_ps2_kb/_0472_ ;
wire \u0_ps2_kb/_0473_ ;
wire \u0_ps2_kb/_0474_ ;
wire \u0_ps2_kb/_0475_ ;
wire \u0_ps2_kb/_0476_ ;
wire \u0_ps2_kb/_0477_ ;
wire \u0_ps2_kb/_0478_ ;
wire \u0_ps2_kb/_0479_ ;
wire \u0_ps2_kb/_0480_ ;
wire \u0_ps2_kb/_0481_ ;
wire \u0_ps2_kb/_0482_ ;
wire \u0_ps2_kb/_0483_ ;
wire \u0_ps2_kb/_0484_ ;
wire \u0_ps2_kb/_0485_ ;
wire \u0_ps2_kb/_0486_ ;
wire \u0_ps2_kb/_0487_ ;
wire \u0_ps2_kb/_0488_ ;
wire \u0_ps2_kb/_0489_ ;
wire \u0_ps2_kb/_0490_ ;
wire \u0_ps2_kb/_0491_ ;
wire \u0_ps2_kb/_0492_ ;
wire \u0_ps2_kb/_0493_ ;
wire \u0_ps2_kb/_0494_ ;
wire \u0_ps2_kb/_0495_ ;
wire \u0_ps2_kb/_0496_ ;
wire \u0_ps2_kb/_0497_ ;
wire \u0_ps2_kb/_0498_ ;
wire \u0_ps2_kb/_0499_ ;
wire \u0_ps2_kb/_0500_ ;
wire \u0_ps2_kb/_0501_ ;
wire \u0_ps2_kb/_0502_ ;
wire \u0_ps2_kb/_0503_ ;
wire \u0_ps2_kb/_0504_ ;
wire \u0_ps2_kb/_0505_ ;
wire \u0_ps2_kb/_0506_ ;
wire \u0_ps2_kb/_0507_ ;
wire \u0_ps2_kb/_0508_ ;
wire \u0_ps2_kb/_0509_ ;
wire \u0_ps2_kb/_0510_ ;
wire \u0_ps2_kb/_0511_ ;
wire \u0_ps2_kb/_0512_ ;
wire \u0_ps2_kb/_0513_ ;
wire \u0_ps2_kb/_0514_ ;
wire \u0_ps2_kb/_0515_ ;
wire \u0_ps2_kb/_0516_ ;
wire \u0_ps2_kb/_0517_ ;
wire \u0_ps2_kb/_0518_ ;
wire \u0_ps2_kb/_0519_ ;
wire \u0_ps2_kb/_0520_ ;
wire \u0_ps2_kb/_0521_ ;
wire \u0_ps2_kb/_0522_ ;
wire \u0_ps2_kb/_0523_ ;
wire \u0_ps2_kb/_0524_ ;
wire \u0_ps2_kb/_0525_ ;
wire \u0_ps2_kb/_0526_ ;
wire \u0_ps2_kb/_0527_ ;
wire \u0_ps2_kb/fifo[0][0] ;
wire \u0_ps2_kb/fifo[0][1] ;
wire \u0_ps2_kb/fifo[0][2] ;
wire \u0_ps2_kb/fifo[0][3] ;
wire \u0_ps2_kb/fifo[0][4] ;
wire \u0_ps2_kb/fifo[0][5] ;
wire \u0_ps2_kb/fifo[0][6] ;
wire \u0_ps2_kb/fifo[0][7] ;
wire \u0_ps2_kb/fifo[1][0] ;
wire \u0_ps2_kb/fifo[1][1] ;
wire \u0_ps2_kb/fifo[1][2] ;
wire \u0_ps2_kb/fifo[1][3] ;
wire \u0_ps2_kb/fifo[1][4] ;
wire \u0_ps2_kb/fifo[1][5] ;
wire \u0_ps2_kb/fifo[1][6] ;
wire \u0_ps2_kb/fifo[1][7] ;
wire \u0_ps2_kb/fifo[2][0] ;
wire \u0_ps2_kb/fifo[2][1] ;
wire \u0_ps2_kb/fifo[2][2] ;
wire \u0_ps2_kb/fifo[2][3] ;
wire \u0_ps2_kb/fifo[2][4] ;
wire \u0_ps2_kb/fifo[2][5] ;
wire \u0_ps2_kb/fifo[2][6] ;
wire \u0_ps2_kb/fifo[2][7] ;
wire \u0_ps2_kb/fifo[3][0] ;
wire \u0_ps2_kb/fifo[3][1] ;
wire \u0_ps2_kb/fifo[3][2] ;
wire \u0_ps2_kb/fifo[3][3] ;
wire \u0_ps2_kb/fifo[3][4] ;
wire \u0_ps2_kb/fifo[3][5] ;
wire \u0_ps2_kb/fifo[3][6] ;
wire \u0_ps2_kb/fifo[3][7] ;
wire \u0_ps2_kb/fifo[4][0] ;
wire \u0_ps2_kb/fifo[4][1] ;
wire \u0_ps2_kb/fifo[4][2] ;
wire \u0_ps2_kb/fifo[4][3] ;
wire \u0_ps2_kb/fifo[4][4] ;
wire \u0_ps2_kb/fifo[4][5] ;
wire \u0_ps2_kb/fifo[4][6] ;
wire \u0_ps2_kb/fifo[4][7] ;
wire \u0_ps2_kb/fifo[5][0] ;
wire \u0_ps2_kb/fifo[5][1] ;
wire \u0_ps2_kb/fifo[5][2] ;
wire \u0_ps2_kb/fifo[5][3] ;
wire \u0_ps2_kb/fifo[5][4] ;
wire \u0_ps2_kb/fifo[5][5] ;
wire \u0_ps2_kb/fifo[5][6] ;
wire \u0_ps2_kb/fifo[5][7] ;
wire \u0_ps2_kb/fifo[6][0] ;
wire \u0_ps2_kb/fifo[6][1] ;
wire \u0_ps2_kb/fifo[6][2] ;
wire \u0_ps2_kb/fifo[6][3] ;
wire \u0_ps2_kb/fifo[6][4] ;
wire \u0_ps2_kb/fifo[6][5] ;
wire \u0_ps2_kb/fifo[6][6] ;
wire \u0_ps2_kb/fifo[6][7] ;
wire \u0_ps2_kb/fifo[7][0] ;
wire \u0_ps2_kb/fifo[7][1] ;
wire \u0_ps2_kb/fifo[7][2] ;
wire \u0_ps2_kb/fifo[7][3] ;
wire \u0_ps2_kb/fifo[7][4] ;
wire \u0_ps2_kb/fifo[7][5] ;
wire \u0_ps2_kb/fifo[7][6] ;
wire \u0_ps2_kb/fifo[7][7] ;
wire \u1_ps2_dsh/_000_ ;
wire \u1_ps2_dsh/_001_ ;
wire \u1_ps2_dsh/_002_ ;
wire \u1_ps2_dsh/_003_ ;
wire \u1_ps2_dsh/_004_ ;
wire \u1_ps2_dsh/_005_ ;
wire \u1_ps2_dsh/_006_ ;
wire \u1_ps2_dsh/_007_ ;
wire \u1_ps2_dsh/_008_ ;
wire \u1_ps2_dsh/_009_ ;
wire \u1_ps2_dsh/_010_ ;
wire \u1_ps2_dsh/_011_ ;
wire \u1_ps2_dsh/_012_ ;
wire \u1_ps2_dsh/_013_ ;
wire \u1_ps2_dsh/_014_ ;
wire \u1_ps2_dsh/_015_ ;
wire \u1_ps2_dsh/_016_ ;
wire \u1_ps2_dsh/_017_ ;
wire \u1_ps2_dsh/_018_ ;
wire \u1_ps2_dsh/_019_ ;
wire \u1_ps2_dsh/_020_ ;
wire \u1_ps2_dsh/_021_ ;
wire \u1_ps2_dsh/_022_ ;
wire \u1_ps2_dsh/_023_ ;
wire \u1_ps2_dsh/_024_ ;
wire \u1_ps2_dsh/_025_ ;
wire \u1_ps2_dsh/_026_ ;
wire \u1_ps2_dsh/_027_ ;
wire \u1_ps2_dsh/_028_ ;
wire \u1_ps2_dsh/_029_ ;
wire \u1_ps2_dsh/_030_ ;
wire \u1_ps2_dsh/_031_ ;
wire \u1_ps2_dsh/_032_ ;
wire \u1_ps2_dsh/_033_ ;
wire \u1_ps2_dsh/_034_ ;
wire \u1_ps2_dsh/_035_ ;
wire \u1_ps2_dsh/_036_ ;
wire \u1_ps2_dsh/_037_ ;
wire \u1_ps2_dsh/_038_ ;
wire \u1_ps2_dsh/_039_ ;
wire \u1_ps2_dsh/_040_ ;
wire \u1_ps2_dsh/_041_ ;
wire \u1_ps2_dsh/_042_ ;
wire \u1_ps2_dsh/_043_ ;
wire \u1_ps2_dsh/_044_ ;
wire \u1_ps2_dsh/_045_ ;
wire \u1_ps2_dsh/_046_ ;
wire \u1_ps2_dsh/_047_ ;
wire \u1_ps2_dsh/_048_ ;
wire \u1_ps2_dsh/_049_ ;
wire \u1_ps2_dsh/_050_ ;
wire \u1_ps2_dsh/_051_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0000_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0001_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0002_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0003_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0004_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0005_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0006_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0007_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0008_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0009_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0010_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0011_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0012_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0013_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0014_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0015_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0016_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0017_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0018_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0019_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0020_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0021_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0022_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0023_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0024_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0025_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0026_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0027_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0028_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0029_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0030_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0031_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0032_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0033_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0034_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0035_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0036_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0037_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0038_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0039_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0040_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0041_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0042_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0043_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0044_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0045_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0046_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0047_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0048_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0049_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0050_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0051_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0052_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0053_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0054_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0055_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0056_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0057_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0058_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0059_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0060_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0061_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0062_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0063_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0064_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0065_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0066_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0067_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0068_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0069_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0070_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0071_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0072_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0073_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0074_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0075_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0076_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0077_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0078_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0079_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0080_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0081_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0082_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0083_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0084_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0085_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0086_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0087_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0088_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0089_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0090_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0091_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0092_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0093_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0094_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0095_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0096_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0097_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0098_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0099_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0100_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0101_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0102_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0103_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0104_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0105_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0106_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0107_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0108_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0109_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0110_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0111_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0112_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0113_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0114_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0115_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0116_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0117_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0118_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0119_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0120_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0121_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0122_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0123_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0124_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0125_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0126_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0127_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0128_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0129_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0130_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0131_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0132_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0133_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0134_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0135_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0136_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0137_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0138_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0139_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0140_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0141_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0142_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0143_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0144_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0145_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0146_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0147_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0148_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0149_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0150_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0151_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0152_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0153_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0154_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0155_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0156_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0157_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0158_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0159_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0160_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0161_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0162_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0163_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0164_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0165_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0166_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0167_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0168_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0169_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0170_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0171_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0172_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0173_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0174_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0175_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0176_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0177_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0178_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0179_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0180_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0181_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0182_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0183_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0184_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0185_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0186_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0187_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0188_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0189_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0190_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0191_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0192_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0193_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0194_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0195_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0196_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0197_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0198_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0199_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0200_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0201_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0202_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0203_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0204_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0205_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0206_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0207_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0208_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0209_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0210_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0211_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0212_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0213_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0214_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0215_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0216_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0217_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0218_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0219_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0220_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0221_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0222_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0223_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0224_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0225_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0226_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0227_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0228_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0229_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0230_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0231_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0232_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0233_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0234_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0235_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0236_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0237_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0238_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0239_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0240_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0241_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0242_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0243_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0244_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0245_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0246_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0247_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0248_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0249_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0250_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0251_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0252_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0253_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0254_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0255_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0256_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0257_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0258_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0259_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0260_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0261_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0262_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0263_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0264_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0265_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0266_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0267_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0268_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0269_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0270_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0271_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0272_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0273_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0274_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0275_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0276_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0277_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0278_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0279_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0280_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0281_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0282_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0283_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0284_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0285_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0286_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0287_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0288_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0289_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0290_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0291_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0292_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0293_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0294_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0295_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0296_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0297_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0298_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0299_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0300_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0301_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0302_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0303_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0304_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0305_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0306_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0307_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0308_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0309_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0310_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0311_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0312_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0313_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0314_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0315_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0316_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0317_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0318_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0319_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0320_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0321_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0322_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0323_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0324_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0325_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0326_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0327_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0328_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0329_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0330_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0331_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0332_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0333_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0334_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0335_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0336_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0337_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0338_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0339_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0340_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0341_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0342_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0343_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0344_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0345_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0346_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0347_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0348_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0349_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0350_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0351_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0352_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0353_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0354_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0355_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0356_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0357_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0358_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0359_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0360_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0361_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0362_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0363_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0364_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0365_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0366_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0367_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0368_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0369_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0370_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0371_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0372_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0373_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0374_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0375_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0376_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0377_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0378_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0379_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0380_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0381_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0382_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0383_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0384_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0385_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0386_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0387_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0388_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0389_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0390_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0391_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0392_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0393_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0394_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0395_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0396_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0397_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0398_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0399_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0400_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0401_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0402_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0403_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0404_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0405_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0406_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0407_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0408_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0409_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0410_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0411_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0412_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0413_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0414_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0415_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0416_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0417_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0418_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0419_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0420_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0421_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0422_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0423_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0424_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0425_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0426_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0427_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0428_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0429_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0430_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0431_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0432_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0433_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0434_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0435_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0436_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0437_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0438_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0439_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0440_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0441_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0442_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0443_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0444_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0445_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0446_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0447_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0448_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0449_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0450_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0451_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0452_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0453_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0454_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0455_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0456_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0457_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0458_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0459_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0460_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0461_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0462_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0463_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0464_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0465_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0466_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0467_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0468_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0469_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0470_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0471_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0472_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0473_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0474_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0475_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0476_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0477_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0478_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0479_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0480_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0481_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0482_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0483_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0484_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0485_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0486_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0487_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0488_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0489_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0490_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0491_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0492_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0493_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0494_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0495_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0496_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0497_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0498_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0499_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0500_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0501_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0502_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0503_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0504_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0505_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0506_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0507_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0508_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0509_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0510_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0511_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0512_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0513_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0514_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0515_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0516_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0517_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0518_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0519_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0520_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0521_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0522_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0523_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0524_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0525_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0526_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0527_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0528_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0529_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0530_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0531_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0532_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0533_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0534_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0535_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0536_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0537_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0538_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0539_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0540_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0541_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0542_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0543_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0544_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0545_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0546_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0547_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0548_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0549_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0550_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0551_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0552_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0553_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0554_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0555_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0556_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0557_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0558_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0559_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0560_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0561_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0562_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0563_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0564_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0565_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0566_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0567_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0568_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0569_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0570_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0571_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0572_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0573_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0574_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0575_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0576_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0577_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0578_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0579_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0580_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0581_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0582_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0583_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0584_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0585_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0586_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0587_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0588_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0589_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0590_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0591_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0592_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0593_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0594_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0595_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0596_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0597_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0598_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0599_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0600_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0601_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0602_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0603_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0604_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0605_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0606_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0607_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0608_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0609_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0610_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0611_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0612_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0613_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0614_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0615_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0616_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0617_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0618_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0619_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0620_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0621_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0622_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0623_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0624_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0625_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0626_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0627_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0628_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0629_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0630_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0631_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0632_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0633_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0634_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0635_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0636_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0637_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0638_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0639_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0640_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0641_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0642_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0643_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0644_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0645_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0646_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0647_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0648_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0649_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0650_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0651_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0652_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0653_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0654_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0655_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0656_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0657_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0658_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0659_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0660_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0661_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0662_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0663_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0664_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0665_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0666_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0667_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0668_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0669_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0670_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0671_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0672_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0673_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0674_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0675_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0676_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0677_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0678_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0679_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0680_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0681_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0682_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0683_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0684_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0685_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0686_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0687_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0688_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0689_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0690_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0691_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0692_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0693_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0694_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0695_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0696_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0697_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0698_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0699_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0700_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0701_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0702_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0703_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0704_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0705_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0706_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0707_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0708_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0709_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0710_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0711_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0712_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0713_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0714_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0715_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0716_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0717_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0718_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0719_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0720_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0721_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0722_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0723_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0724_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0725_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0726_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0727_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0728_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0729_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0730_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0731_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0732_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0733_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0734_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0735_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0736_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0737_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0738_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0739_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0740_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0741_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0742_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0743_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0744_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0745_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0746_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0747_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0748_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0749_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0750_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0751_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0752_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0753_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0754_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0755_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0756_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0757_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0758_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0759_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0760_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0761_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0762_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0763_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0764_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0765_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0766_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0767_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0768_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0769_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0770_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0771_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0772_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0773_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0774_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0775_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0776_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0777_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0778_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0779_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0780_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0781_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0782_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0783_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0784_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0785_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0786_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0787_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0788_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0789_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0790_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0791_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0792_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0793_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0794_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0795_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0796_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0797_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0798_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0799_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0800_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0801_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0802_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0803_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0804_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0805_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0806_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0807_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0808_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0809_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0810_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0811_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0812_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0813_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0814_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0815_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0816_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0817_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0818_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0819_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0820_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0821_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0822_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0823_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0824_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0825_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0826_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0827_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0828_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0829_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0830_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0831_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0832_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0833_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0834_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0835_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0836_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0837_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0838_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0839_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0840_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0841_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0842_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0843_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0844_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0845_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0846_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0847_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0848_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0849_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0850_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0851_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0852_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0853_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0854_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0855_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0856_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0857_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0858_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0859_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0860_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0861_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0862_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0863_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0864_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0865_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0866_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0867_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0868_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0869_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0870_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0871_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0872_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0873_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0874_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0875_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0876_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0877_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0878_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0879_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0880_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0881_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0882_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0883_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0884_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0885_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0886_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0887_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0888_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0889_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0890_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0891_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0892_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0893_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0894_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0895_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0896_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0897_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0898_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0899_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0900_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0901_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0902_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0903_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0904_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0905_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0906_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0907_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0908_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0909_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0910_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0911_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0912_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0913_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0914_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0915_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0916_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0917_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0918_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0919_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0920_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0921_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0922_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0923_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0924_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0925_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0926_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0927_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0928_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0929_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0930_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0931_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0932_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0933_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0934_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0935_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0936_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0937_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0938_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0939_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0940_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0941_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0942_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0943_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0944_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0945_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0946_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0947_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0948_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0949_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0950_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0951_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0952_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0953_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0954_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0955_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0956_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0957_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0958_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0959_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0960_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0961_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0962_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0963_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0964_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0965_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0966_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0967_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0968_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0969_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0970_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0971_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0972_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0973_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0974_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0975_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0976_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0977_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0978_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0979_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0980_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0981_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0982_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0983_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0984_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0985_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0986_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0987_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0988_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0989_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0990_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0991_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0992_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0993_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0994_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0995_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0996_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0997_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0998_ ;
wire \u1_ps2_dsh/key_ascii/i0/_0999_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1000_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1001_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1002_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1003_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1004_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1005_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1006_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1007_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1008_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1009_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1010_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1011_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1012_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1013_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1014_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1015_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1016_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1017_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1018_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1019_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1020_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1021_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1022_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1023_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1024_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1025_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1026_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1027_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1028_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1029_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1030_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1031_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1032_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1033_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1034_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1035_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1036_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1037_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1038_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1039_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1040_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1041_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1042_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1043_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1044_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1045_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1046_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1047_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1048_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1049_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1050_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1051_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1052_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1053_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1054_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1055_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1056_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1057_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1058_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1059_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1060_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1061_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1062_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1063_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1064_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1065_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1066_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1067_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1068_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1069_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1070_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1071_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1072_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1073_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1074_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1075_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1076_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1077_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1078_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1079_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1080_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1081_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1082_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1083_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1084_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1085_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1086_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1087_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1088_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1089_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1090_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1091_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1092_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1093_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1094_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1095_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1096_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1097_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1098_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1099_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1100_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1101_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1102_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1103_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1104_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1105_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1106_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1107_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1108_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1109_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1110_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1111_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1112_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1113_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1114_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1115_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1116_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1117_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1118_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1119_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1120_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1121_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1122_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1123_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1124_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1125_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1126_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1127_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1128_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1129_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1130_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1131_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1132_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1133_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1134_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1135_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1136_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1137_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1138_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1139_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1140_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1141_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1142_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1143_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1144_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1145_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1146_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1147_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1148_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1149_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1150_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1151_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1152_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1153_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1154_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1155_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1156_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1157_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1158_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1159_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1160_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1161_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1162_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1163_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1164_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1165_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1166_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1167_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1168_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1169_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1170_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1171_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1172_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1173_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1174_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1175_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1176_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1177_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1178_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1179_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1180_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1181_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1182_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1183_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1184_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1185_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1186_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1187_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1188_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1189_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1190_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1191_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1192_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1193_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1194_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1195_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1196_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1197_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1198_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1199_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1200_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1201_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1202_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1203_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1204_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1205_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1206_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1207_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1208_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1209_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1210_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1211_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1212_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1213_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1214_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1215_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1216_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1217_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1218_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1219_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1220_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1221_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1222_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1223_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1224_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1225_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1226_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1227_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1228_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1229_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1230_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1231_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1232_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1233_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1234_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1235_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1236_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1237_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1238_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1239_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1240_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1241_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1242_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1243_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1244_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1245_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1246_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1247_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1248_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1249_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1250_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1251_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1252_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1253_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1254_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1255_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1256_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1257_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1258_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1259_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1260_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1261_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1262_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1263_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1264_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1265_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1266_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1267_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1268_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1269_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1270_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1271_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1272_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1273_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1274_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1275_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1276_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1277_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1278_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1279_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1280_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1281_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1282_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1283_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1284_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1285_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1286_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1287_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1288_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1289_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1290_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1291_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1292_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1293_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1294_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1295_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1296_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1297_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1298_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1299_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1300_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1301_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1302_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1303_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1304_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1305_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1306_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1307_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1308_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1309_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1310_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1311_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1312_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1313_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1314_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1315_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1316_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1317_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1318_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1319_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1320_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1321_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1322_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1323_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1324_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1325_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1326_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1327_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1328_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1329_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1330_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1331_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1332_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1333_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1334_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1335_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1336_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1337_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1338_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1339_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1340_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1341_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1342_ ;
wire \u1_ps2_dsh/key_ascii/i0/_1343_ ;
wire \u2_ps2_cer/_000_ ;
wire \u2_ps2_cer/_001_ ;
wire \u2_ps2_cer/_002_ ;
wire \u2_ps2_cer/_003_ ;
wire \u2_ps2_cer/_004_ ;
wire \u2_ps2_cer/_005_ ;
wire \u2_ps2_cer/_006_ ;
wire \u2_ps2_cer/_007_ ;
wire \u2_ps2_cer/_008_ ;
wire \u2_ps2_cer/_009_ ;
wire \u2_ps2_cer/_010_ ;
wire \u2_ps2_cer/_011_ ;
wire \u2_ps2_cer/_012_ ;
wire \u2_ps2_cer/_013_ ;
wire \u2_ps2_cer/_014_ ;
wire \u2_ps2_cer/_015_ ;
wire \u2_ps2_cer/_016_ ;
wire \u2_ps2_cer/_017_ ;
wire \u2_ps2_cer/_018_ ;
wire \u2_ps2_cer/_019_ ;
wire \u2_ps2_cer/_020_ ;
wire \u2_ps2_cer/_021_ ;
wire \u2_ps2_cer/_022_ ;
wire \u2_ps2_cer/_023_ ;
wire \u2_ps2_cer/_024_ ;
wire \u2_ps2_cer/_025_ ;
wire \u2_ps2_cer/_026_ ;
wire \u2_ps2_cer/_027_ ;
wire \u2_ps2_cer/_028_ ;
wire \u2_ps2_cer/_029_ ;
wire \u2_ps2_cer/_030_ ;
wire \u2_ps2_cer/_031_ ;
wire \u2_ps2_cer/_032_ ;
wire \u2_ps2_cer/_033_ ;
wire \u2_ps2_cer/_034_ ;
wire \u2_ps2_cer/_035_ ;
wire \u2_ps2_cer/_036_ ;
wire \u2_ps2_cer/_037_ ;
wire \u2_ps2_cer/_038_ ;
wire \u2_ps2_cer/_039_ ;
wire \u2_ps2_cer/_040_ ;
wire \u2_ps2_cer/_041_ ;
wire \u2_ps2_cer/_042_ ;
wire \u2_ps2_cer/_043_ ;
wire \u2_ps2_cer/_044_ ;
wire \u2_ps2_cer/_045_ ;
wire \u2_ps2_cer/_046_ ;
wire \u2_ps2_cer/_047_ ;
wire \u2_ps2_cer/_048_ ;
wire \u2_ps2_cer/_049_ ;
wire \u2_ps2_cer/_050_ ;
wire \u2_ps2_cer/_051_ ;
wire \u2_ps2_cer/_052_ ;
wire \u2_ps2_cer/_053_ ;
wire \u2_ps2_cer/_054_ ;
wire \u2_ps2_cer/_055_ ;
wire \u2_ps2_cer/_056_ ;
wire \u2_ps2_cer/_057_ ;
wire \u2_ps2_cer/_058_ ;
wire \u2_ps2_cer/_059_ ;
wire \u2_ps2_cer/_060_ ;
wire \u2_ps2_cer/_061_ ;
wire \u2_ps2_cer/_062_ ;
wire \u2_ps2_cer/_063_ ;
wire \u2_ps2_cer/_064_ ;
wire \u2_ps2_cer/_065_ ;
wire \u2_ps2_cer/_066_ ;
wire \u2_ps2_cer/counted ;
wire \u3_seg_h_0/_00_ ;
wire \u3_seg_h_0/_01_ ;
wire \u3_seg_h_0/_02_ ;
wire \u3_seg_h_0/_03_ ;
wire \u3_seg_h_0/_04_ ;
wire \u3_seg_h_0/_05_ ;
wire \u3_seg_h_0/_06_ ;
wire \u3_seg_h_0/_07_ ;
wire \u3_seg_h_0/_08_ ;
wire \u3_seg_h_0/_09_ ;
wire \u3_seg_h_0/_10_ ;
wire \u3_seg_h_0/_11_ ;
wire \u3_seg_h_0/_12_ ;
wire \u3_seg_h_0/_13_ ;
wire \u3_seg_h_0/_14_ ;
wire \u3_seg_h_0/_15_ ;
wire \u3_seg_h_0/_16_ ;
wire \u3_seg_h_0/_17_ ;
wire \u3_seg_h_0/_18_ ;
wire \u3_seg_h_0/_19_ ;
wire \u3_seg_h_0/_20_ ;
wire \u3_seg_h_0/_21_ ;
wire \u3_seg_h_0/_22_ ;
wire \u3_seg_h_0/_23_ ;
wire \u3_seg_h_0/_24_ ;
wire \u3_seg_h_0/_25_ ;
wire \u3_seg_h_0/_26_ ;
wire \u3_seg_h_0/_27_ ;
wire \u3_seg_h_0/_28_ ;
wire \u3_seg_h_0/_29_ ;
wire \u3_seg_h_0/_30_ ;
wire \u3_seg_h_0/_31_ ;
wire \u3_seg_h_0/_32_ ;
wire \u3_seg_h_0/_33_ ;
wire \u3_seg_h_0/_34_ ;
wire \u3_seg_h_0/_35_ ;
wire \u3_seg_h_0/_36_ ;
wire \u3_seg_h_0/_37_ ;
wire \u3_seg_h_0/_38_ ;
wire \u3_seg_h_0/_39_ ;
wire \u3_seg_h_0/_40_ ;
wire \u3_seg_h_0/_41_ ;
wire \u3_seg_h_0/_42_ ;
wire \u4_seg_h_1/_00_ ;
wire \u4_seg_h_1/_01_ ;
wire \u4_seg_h_1/_02_ ;
wire \u4_seg_h_1/_03_ ;
wire \u4_seg_h_1/_04_ ;
wire \u4_seg_h_1/_05_ ;
wire \u4_seg_h_1/_06_ ;
wire \u4_seg_h_1/_07_ ;
wire \u4_seg_h_1/_08_ ;
wire \u4_seg_h_1/_09_ ;
wire \u4_seg_h_1/_10_ ;
wire \u4_seg_h_1/_11_ ;
wire \u4_seg_h_1/_12_ ;
wire \u4_seg_h_1/_13_ ;
wire \u4_seg_h_1/_14_ ;
wire \u4_seg_h_1/_15_ ;
wire \u4_seg_h_1/_16_ ;
wire \u4_seg_h_1/_17_ ;
wire \u4_seg_h_1/_18_ ;
wire \u4_seg_h_1/_19_ ;
wire \u4_seg_h_1/_20_ ;
wire \u4_seg_h_1/_21_ ;
wire \u4_seg_h_1/_22_ ;
wire \u4_seg_h_1/_23_ ;
wire \u4_seg_h_1/_24_ ;
wire \u4_seg_h_1/_25_ ;
wire \u4_seg_h_1/_26_ ;
wire \u4_seg_h_1/_27_ ;
wire \u4_seg_h_1/_28_ ;
wire \u4_seg_h_1/_29_ ;
wire \u4_seg_h_1/_30_ ;
wire \u4_seg_h_1/_31_ ;
wire \u4_seg_h_1/_32_ ;
wire \u4_seg_h_1/_33_ ;
wire \u4_seg_h_1/_34_ ;
wire \u4_seg_h_1/_35_ ;
wire \u4_seg_h_1/_36_ ;
wire \u4_seg_h_1/_37_ ;
wire \u4_seg_h_1/_38_ ;
wire \u4_seg_h_1/_39_ ;
wire \u4_seg_h_1/_40_ ;
wire \u4_seg_h_1/_41_ ;
wire \u4_seg_h_1/_42_ ;
wire \u5_seg_h_2/_00_ ;
wire \u5_seg_h_2/_01_ ;
wire \u5_seg_h_2/_02_ ;
wire \u5_seg_h_2/_03_ ;
wire \u5_seg_h_2/_04_ ;
wire \u5_seg_h_2/_05_ ;
wire \u5_seg_h_2/_06_ ;
wire \u5_seg_h_2/_07_ ;
wire \u5_seg_h_2/_08_ ;
wire \u5_seg_h_2/_09_ ;
wire \u5_seg_h_2/_10_ ;
wire \u5_seg_h_2/_11_ ;
wire \u5_seg_h_2/_12_ ;
wire \u5_seg_h_2/_13_ ;
wire \u5_seg_h_2/_14_ ;
wire \u5_seg_h_2/_15_ ;
wire \u5_seg_h_2/_16_ ;
wire \u5_seg_h_2/_17_ ;
wire \u5_seg_h_2/_18_ ;
wire \u5_seg_h_2/_19_ ;
wire \u5_seg_h_2/_20_ ;
wire \u5_seg_h_2/_21_ ;
wire \u5_seg_h_2/_22_ ;
wire \u5_seg_h_2/_23_ ;
wire \u5_seg_h_2/_24_ ;
wire \u5_seg_h_2/_25_ ;
wire \u5_seg_h_2/_26_ ;
wire \u5_seg_h_2/_27_ ;
wire \u5_seg_h_2/_28_ ;
wire \u5_seg_h_2/_29_ ;
wire \u5_seg_h_2/_30_ ;
wire \u5_seg_h_2/_31_ ;
wire \u5_seg_h_2/_32_ ;
wire \u5_seg_h_2/_33_ ;
wire \u5_seg_h_2/_34_ ;
wire \u5_seg_h_2/_35_ ;
wire \u5_seg_h_2/_36_ ;
wire \u5_seg_h_2/_37_ ;
wire \u5_seg_h_2/_38_ ;
wire \u5_seg_h_2/_39_ ;
wire \u5_seg_h_2/_40_ ;
wire \u5_seg_h_2/_41_ ;
wire \u5_seg_h_2/_42_ ;
wire \u6_seg_h_3/_00_ ;
wire \u6_seg_h_3/_01_ ;
wire \u6_seg_h_3/_02_ ;
wire \u6_seg_h_3/_03_ ;
wire \u6_seg_h_3/_04_ ;
wire \u6_seg_h_3/_05_ ;
wire \u6_seg_h_3/_06_ ;
wire \u6_seg_h_3/_07_ ;
wire \u6_seg_h_3/_08_ ;
wire \u6_seg_h_3/_09_ ;
wire \u6_seg_h_3/_10_ ;
wire \u6_seg_h_3/_11_ ;
wire \u6_seg_h_3/_12_ ;
wire \u6_seg_h_3/_13_ ;
wire \u6_seg_h_3/_14_ ;
wire \u6_seg_h_3/_15_ ;
wire \u6_seg_h_3/_16_ ;
wire \u6_seg_h_3/_17_ ;
wire \u6_seg_h_3/_18_ ;
wire \u6_seg_h_3/_19_ ;
wire \u6_seg_h_3/_20_ ;
wire \u6_seg_h_3/_21_ ;
wire \u6_seg_h_3/_22_ ;
wire \u6_seg_h_3/_23_ ;
wire \u6_seg_h_3/_24_ ;
wire \u6_seg_h_3/_25_ ;
wire \u6_seg_h_3/_26_ ;
wire \u6_seg_h_3/_27_ ;
wire \u6_seg_h_3/_28_ ;
wire \u6_seg_h_3/_29_ ;
wire \u6_seg_h_3/_30_ ;
wire \u6_seg_h_3/_31_ ;
wire \u6_seg_h_3/_32_ ;
wire \u6_seg_h_3/_33_ ;
wire \u6_seg_h_3/_34_ ;
wire \u6_seg_h_3/_35_ ;
wire \u6_seg_h_3/_36_ ;
wire \u6_seg_h_3/_37_ ;
wire \u6_seg_h_3/_38_ ;
wire \u6_seg_h_3/_39_ ;
wire \u6_seg_h_3/_40_ ;
wire \u6_seg_h_3/_41_ ;
wire \u6_seg_h_3/_42_ ;
wire \u7_seg_h_4/_00_ ;
wire \u7_seg_h_4/_01_ ;
wire \u7_seg_h_4/_02_ ;
wire \u7_seg_h_4/_03_ ;
wire \u7_seg_h_4/_04_ ;
wire \u7_seg_h_4/_05_ ;
wire \u7_seg_h_4/_06_ ;
wire \u7_seg_h_4/_07_ ;
wire \u7_seg_h_4/_08_ ;
wire \u7_seg_h_4/_09_ ;
wire \u7_seg_h_4/_10_ ;
wire \u7_seg_h_4/_11_ ;
wire \u7_seg_h_4/_12_ ;
wire \u7_seg_h_4/_13_ ;
wire \u7_seg_h_4/_14_ ;
wire \u7_seg_h_4/_15_ ;
wire \u7_seg_h_4/_16_ ;
wire \u7_seg_h_4/_17_ ;
wire \u7_seg_h_4/_18_ ;
wire \u7_seg_h_4/_19_ ;
wire \u7_seg_h_4/_20_ ;
wire \u7_seg_h_4/_21_ ;
wire \u7_seg_h_4/_22_ ;
wire \u7_seg_h_4/_23_ ;
wire \u7_seg_h_4/_24_ ;
wire \u7_seg_h_4/_25_ ;
wire \u7_seg_h_4/_26_ ;
wire \u7_seg_h_4/_27_ ;
wire \u7_seg_h_4/_28_ ;
wire \u7_seg_h_4/_29_ ;
wire \u7_seg_h_4/_30_ ;
wire \u7_seg_h_4/_31_ ;
wire \u7_seg_h_4/_32_ ;
wire \u7_seg_h_4/_33_ ;
wire \u7_seg_h_4/_34_ ;
wire \u7_seg_h_4/_35_ ;
wire \u7_seg_h_4/_36_ ;
wire \u7_seg_h_4/_37_ ;
wire \u7_seg_h_4/_38_ ;
wire \u7_seg_h_4/_39_ ;
wire \u7_seg_h_4/_40_ ;
wire \u7_seg_h_4/_41_ ;
wire \u7_seg_h_4/_42_ ;
wire \u8_seg_h_5/_00_ ;
wire \u8_seg_h_5/_01_ ;
wire \u8_seg_h_5/_02_ ;
wire \u8_seg_h_5/_03_ ;
wire \u8_seg_h_5/_04_ ;
wire \u8_seg_h_5/_05_ ;
wire \u8_seg_h_5/_06_ ;
wire \u8_seg_h_5/_07_ ;
wire \u8_seg_h_5/_08_ ;
wire \u8_seg_h_5/_09_ ;
wire \u8_seg_h_5/_10_ ;
wire \u8_seg_h_5/_11_ ;
wire \u8_seg_h_5/_12_ ;
wire \u8_seg_h_5/_13_ ;
wire \u8_seg_h_5/_14_ ;
wire \u8_seg_h_5/_15_ ;
wire \u8_seg_h_5/_16_ ;
wire \u8_seg_h_5/_17_ ;
wire \u8_seg_h_5/_18_ ;
wire \u8_seg_h_5/_19_ ;
wire \u8_seg_h_5/_20_ ;
wire \u8_seg_h_5/_21_ ;
wire \u8_seg_h_5/_22_ ;
wire \u8_seg_h_5/_23_ ;
wire \u8_seg_h_5/_24_ ;
wire \u8_seg_h_5/_25_ ;
wire \u8_seg_h_5/_26_ ;
wire \u8_seg_h_5/_27_ ;
wire \u8_seg_h_5/_28_ ;
wire \u8_seg_h_5/_29_ ;
wire \u8_seg_h_5/_30_ ;
wire \u8_seg_h_5/_31_ ;
wire \u8_seg_h_5/_32_ ;
wire \u8_seg_h_5/_33_ ;
wire \u8_seg_h_5/_34_ ;
wire \u8_seg_h_5/_35_ ;
wire \u8_seg_h_5/_36_ ;
wire \u8_seg_h_5/_37_ ;
wire \u8_seg_h_5/_38_ ;
wire \u8_seg_h_5/_39_ ;
wire \u8_seg_h_5/_40_ ;
wire \u8_seg_h_5/_41_ ;
wire \u8_seg_h_5/_42_ ;
wire clk ;
wire clrn ;
wire ps2_data ;
wire overflow ;
wire ps2_clk ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire [7:0] ascii ;
wire [7:0] data ;
wire [7:0] data_d1 ;
wire [3:0] high_tens ;
wire [3:0] high_units ;
wire [7:0] key_ascii_display ;
wire [7:0] key_scan_display ;
wire [9:0] \u0_ps2_kb/buffer ;
wire [3:0] \u0_ps2_kb/count ;
wire [2:0] \u0_ps2_kb/ps2_clk_sync ;
wire [2:0] \u0_ps2_kb/r_ptr ;
wire [2:0] \u0_ps2_kb/w_ptr ;
wire [7:0] \u1_ps2_dsh/ascii_result ;
wire [7:0] seg_out_2 ;
wire [7:0] seg_out_3 ;
wire [7:0] seg_out_0 ;
wire [7:0] seg_out_1 ;
wire [7:0] seg_out_4 ;
wire [7:0] seg_out_5 ;


INV_X32 _133_ ( .A(_103_ ), .ZN(_098_ ) );
NOR3_X1 _134_ ( .A1(_098_ ), .A2(_104_ ), .A3(_087_ ), .ZN(_053_ ) );
NOR2_X4 _135_ ( .A1(_098_ ), .A2(_104_ ), .ZN(_099_ ) );
BUF_X4 _136_ ( .A(_099_ ), .Z(_100_ ) );
MUX2_X1 _137_ ( .A(_070_ ), .B(_062_ ), .S(_100_ ), .Z(_027_ ) );
MUX2_X1 _138_ ( .A(_071_ ), .B(_063_ ), .S(_100_ ), .Z(_028_ ) );
MUX2_X1 _139_ ( .A(_072_ ), .B(_064_ ), .S(_100_ ), .Z(_029_ ) );
MUX2_X1 _140_ ( .A(_073_ ), .B(_065_ ), .S(_100_ ), .Z(_030_ ) );
MUX2_X1 _141_ ( .A(_074_ ), .B(_066_ ), .S(_100_ ), .Z(_031_ ) );
MUX2_X1 _142_ ( .A(_075_ ), .B(_067_ ), .S(_100_ ), .Z(_032_ ) );
MUX2_X1 _143_ ( .A(_076_ ), .B(_068_ ), .S(_100_ ), .Z(_033_ ) );
MUX2_X1 _144_ ( .A(_077_ ), .B(_069_ ), .S(_100_ ), .Z(_034_ ) );
MUX2_X1 _145_ ( .A(_079_ ), .B(_054_ ), .S(_100_ ), .Z(_036_ ) );
BUF_X4 _146_ ( .A(_099_ ), .Z(_101_ ) );
MUX2_X1 _147_ ( .A(_080_ ), .B(_055_ ), .S(_101_ ), .Z(_037_ ) );
MUX2_X1 _148_ ( .A(_081_ ), .B(_056_ ), .S(_101_ ), .Z(_038_ ) );
MUX2_X1 _149_ ( .A(_082_ ), .B(_057_ ), .S(_101_ ), .Z(_039_ ) );
MUX2_X1 _150_ ( .A(_083_ ), .B(_058_ ), .S(_101_ ), .Z(_040_ ) );
MUX2_X1 _151_ ( .A(_084_ ), .B(_059_ ), .S(_101_ ), .Z(_041_ ) );
MUX2_X1 _152_ ( .A(_085_ ), .B(_060_ ), .S(_101_ ), .Z(_042_ ) );
MUX2_X1 _153_ ( .A(_086_ ), .B(_061_ ), .S(_101_ ), .Z(_043_ ) );
MUX2_X1 _154_ ( .A(_088_ ), .B(_062_ ), .S(_101_ ), .Z(_044_ ) );
MUX2_X1 _155_ ( .A(_089_ ), .B(_063_ ), .S(_101_ ), .Z(_045_ ) );
MUX2_X1 _156_ ( .A(_090_ ), .B(_064_ ), .S(_101_ ), .Z(_046_ ) );
MUX2_X1 _157_ ( .A(_091_ ), .B(_065_ ), .S(_099_ ), .Z(_047_ ) );
MUX2_X1 _158_ ( .A(_092_ ), .B(_066_ ), .S(_099_ ), .Z(_048_ ) );
MUX2_X1 _159_ ( .A(_093_ ), .B(_067_ ), .S(_099_ ), .Z(_049_ ) );
MUX2_X1 _160_ ( .A(_094_ ), .B(_068_ ), .S(_099_ ), .Z(_050_ ) );
MUX2_X1 _161_ ( .A(_095_ ), .B(_069_ ), .S(_099_ ), .Z(_051_ ) );
INV_X1 _162_ ( .A(_102_ ), .ZN(_096_ ) );
AOI21_X1 _163_ ( .A(_100_ ), .B1(_087_ ), .B2(_096_ ), .ZN(_052_ ) );
INV_X1 _164_ ( .A(_078_ ), .ZN(_097_ ) );
OAI22_X1 _165_ ( .A1(_098_ ), .A2(_104_ ), .B1(_097_ ), .B2(_087_ ), .ZN(_035_ ) );
LOGIC1_X1 _166_ ( .Z(_132_ ) );
BUF_X1 _167_ ( .A(ready ), .Z(_103_ ) );
BUF_X1 _168_ ( .A(ready_d1 ), .Z(_104_ ) );
BUF_X1 _169_ ( .A(key_release ), .Z(_087_ ) );
BUF_X1 _170_ ( .A(_053_ ), .Z(_026_ ) );
BUF_X1 _171_ ( .A(\data [0] ), .Z(_062_ ) );
BUF_X1 _172_ ( .A(\data_d1 [0] ), .Z(_070_ ) );
BUF_X1 _173_ ( .A(_027_ ), .Z(_000_ ) );
BUF_X1 _174_ ( .A(\data [1] ), .Z(_063_ ) );
BUF_X1 _175_ ( .A(\data_d1 [1] ), .Z(_071_ ) );
BUF_X1 _176_ ( .A(_028_ ), .Z(_001_ ) );
BUF_X1 _177_ ( .A(\data [2] ), .Z(_064_ ) );
BUF_X1 _178_ ( .A(\data_d1 [2] ), .Z(_072_ ) );
BUF_X1 _179_ ( .A(_029_ ), .Z(_002_ ) );
BUF_X1 _180_ ( .A(\data [3] ), .Z(_065_ ) );
BUF_X1 _181_ ( .A(\data_d1 [3] ), .Z(_073_ ) );
BUF_X1 _182_ ( .A(_030_ ), .Z(_003_ ) );
BUF_X1 _183_ ( .A(\data [4] ), .Z(_066_ ) );
BUF_X1 _184_ ( .A(\data_d1 [4] ), .Z(_074_ ) );
BUF_X1 _185_ ( .A(_031_ ), .Z(_004_ ) );
BUF_X1 _186_ ( .A(\data [5] ), .Z(_067_ ) );
BUF_X1 _187_ ( .A(\data_d1 [5] ), .Z(_075_ ) );
BUF_X1 _188_ ( .A(_032_ ), .Z(_005_ ) );
BUF_X1 _189_ ( .A(\data [6] ), .Z(_068_ ) );
BUF_X1 _190_ ( .A(\data_d1 [6] ), .Z(_076_ ) );
BUF_X1 _191_ ( .A(_033_ ), .Z(_006_ ) );
BUF_X1 _192_ ( .A(\data [7] ), .Z(_069_ ) );
BUF_X1 _193_ ( .A(\data_d1 [7] ), .Z(_077_ ) );
BUF_X1 _194_ ( .A(_034_ ), .Z(_007_ ) );
BUF_X1 _195_ ( .A(\ascii [0] ), .Z(_054_ ) );
BUF_X1 _196_ ( .A(\key_ascii_display [0] ), .Z(_079_ ) );
BUF_X1 _197_ ( .A(_036_ ), .Z(_009_ ) );
BUF_X1 _198_ ( .A(\ascii [1] ), .Z(_055_ ) );
BUF_X1 _199_ ( .A(\key_ascii_display [1] ), .Z(_080_ ) );
BUF_X1 _200_ ( .A(_037_ ), .Z(_010_ ) );
BUF_X1 _201_ ( .A(\ascii [2] ), .Z(_056_ ) );
BUF_X1 _202_ ( .A(\key_ascii_display [2] ), .Z(_081_ ) );
BUF_X1 _203_ ( .A(_038_ ), .Z(_011_ ) );
BUF_X1 _204_ ( .A(\ascii [3] ), .Z(_057_ ) );
BUF_X1 _205_ ( .A(\key_ascii_display [3] ), .Z(_082_ ) );
BUF_X1 _206_ ( .A(_039_ ), .Z(_012_ ) );
BUF_X1 _207_ ( .A(\ascii [4] ), .Z(_058_ ) );
BUF_X1 _208_ ( .A(\key_ascii_display [4] ), .Z(_083_ ) );
BUF_X1 _209_ ( .A(_040_ ), .Z(_013_ ) );
BUF_X1 _210_ ( .A(\ascii [5] ), .Z(_059_ ) );
BUF_X1 _211_ ( .A(\key_ascii_display [5] ), .Z(_084_ ) );
BUF_X1 _212_ ( .A(_041_ ), .Z(_014_ ) );
BUF_X1 _213_ ( .A(\ascii [6] ), .Z(_060_ ) );
BUF_X1 _214_ ( .A(\key_ascii_display [6] ), .Z(_085_ ) );
BUF_X1 _215_ ( .A(_042_ ), .Z(_015_ ) );
BUF_X1 _216_ ( .A(\ascii [7] ), .Z(_061_ ) );
BUF_X1 _217_ ( .A(\key_ascii_display [7] ), .Z(_086_ ) );
BUF_X1 _218_ ( .A(_043_ ), .Z(_016_ ) );
BUF_X1 _219_ ( .A(\key_scan_display [0] ), .Z(_088_ ) );
BUF_X1 _220_ ( .A(_044_ ), .Z(_017_ ) );
BUF_X1 _221_ ( .A(\key_scan_display [1] ), .Z(_089_ ) );
BUF_X1 _222_ ( .A(_045_ ), .Z(_018_ ) );
BUF_X1 _223_ ( .A(\key_scan_display [2] ), .Z(_090_ ) );
BUF_X1 _224_ ( .A(_046_ ), .Z(_019_ ) );
BUF_X1 _225_ ( .A(\key_scan_display [3] ), .Z(_091_ ) );
BUF_X1 _226_ ( .A(_047_ ), .Z(_020_ ) );
BUF_X1 _227_ ( .A(\key_scan_display [4] ), .Z(_092_ ) );
BUF_X1 _228_ ( .A(_048_ ), .Z(_021_ ) );
BUF_X1 _229_ ( .A(\key_scan_display [5] ), .Z(_093_ ) );
BUF_X1 _230_ ( .A(_049_ ), .Z(_022_ ) );
BUF_X1 _231_ ( .A(\key_scan_display [6] ), .Z(_094_ ) );
BUF_X1 _232_ ( .A(_050_ ), .Z(_023_ ) );
BUF_X1 _233_ ( .A(\key_scan_display [7] ), .Z(_095_ ) );
BUF_X1 _234_ ( .A(_051_ ), .Z(_024_ ) );
BUF_X1 _235_ ( .A(nextdata_n ), .Z(_102_ ) );
BUF_X1 _236_ ( .A(_052_ ), .Z(_025_ ) );
BUF_X1 _237_ ( .A(en ), .Z(_078_ ) );
BUF_X1 _238_ ( .A(_035_ ), .Z(_008_ ) );
DFFS_X1 _239_ ( .D(_025_ ), .SN(fanout_net_28 ), .CK(clk ), .Q(nextdata_n ), .QN(_105_ ) );
DFFR_X1 _240_ ( .D(_000_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [0] ), .QN(_106_ ) );
DFFR_X1 _241_ ( .D(_001_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [1] ), .QN(_107_ ) );
DFFR_X1 _242_ ( .D(_002_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [2] ), .QN(_108_ ) );
DFFR_X1 _243_ ( .D(_003_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [3] ), .QN(_109_ ) );
DFFR_X1 _244_ ( .D(_004_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [4] ), .QN(_110_ ) );
DFFR_X1 _245_ ( .D(_005_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [5] ), .QN(_111_ ) );
DFFR_X1 _246_ ( .D(_006_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [6] ), .QN(_112_ ) );
DFFR_X1 _247_ ( .D(_007_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\data_d1 [7] ), .QN(_113_ ) );
DFFR_X1 _248_ ( .D(_017_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [0] ), .QN(_114_ ) );
DFFR_X1 _249_ ( .D(_018_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [1] ), .QN(_115_ ) );
DFFR_X1 _250_ ( .D(_019_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [2] ), .QN(_116_ ) );
DFFR_X1 _251_ ( .D(_020_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [3] ), .QN(_117_ ) );
DFFR_X1 _252_ ( .D(_021_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [4] ), .QN(_118_ ) );
DFFR_X1 _253_ ( .D(_022_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [5] ), .QN(_119_ ) );
DFFR_X1 _254_ ( .D(_023_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [6] ), .QN(_120_ ) );
DFFR_X1 _255_ ( .D(_024_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_scan_display [7] ), .QN(_121_ ) );
DFFR_X1 _256_ ( .D(_009_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [0] ), .QN(_122_ ) );
DFFR_X1 _257_ ( .D(_010_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [1] ), .QN(_123_ ) );
DFFR_X1 _258_ ( .D(_011_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [2] ), .QN(_124_ ) );
DFFR_X1 _259_ ( .D(_012_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [3] ), .QN(_125_ ) );
DFFR_X1 _260_ ( .D(_013_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [4] ), .QN(_126_ ) );
DFFR_X1 _261_ ( .D(_014_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [5] ), .QN(_127_ ) );
DFFR_X1 _262_ ( .D(_015_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [6] ), .QN(_128_ ) );
DFFR_X1 _263_ ( .D(_016_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\key_ascii_display [7] ), .QN(_129_ ) );
DFFR_X1 _264_ ( .D(_008_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(en ), .QN(_130_ ) );
DFFR_X1 _265_ ( .D(ready ), .RN(fanout_net_28 ), .CK(clk ), .Q(ready_d1 ), .QN(_131_ ) );
INV_X1 \u0_ps2_kb/_0528_ ( .A(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0279_ ) );
NOR2_X1 \u0_ps2_kb/_0529_ ( .A1(\u0_ps2_kb/_0279_ ), .A2(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0280_ ) );
INV_X1 \u0_ps2_kb/_0530_ ( .A(\u0_ps2_kb/_0206_ ), .ZN(\u0_ps2_kb/_0281_ ) );
AND3_X1 \u0_ps2_kb/_0531_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0205_ ), .A3(\u0_ps2_kb/_0281_ ), .ZN(\u0_ps2_kb/_0282_ ) );
INV_X1 \u0_ps2_kb/_0532_ ( .A(\u0_ps2_kb/_0440_ ), .ZN(\u0_ps2_kb/_0283_ ) );
NOR2_X1 \u0_ps2_kb/_0533_ ( .A1(\u0_ps2_kb/_0283_ ), .A2(\u0_ps2_kb/_0439_ ), .ZN(\u0_ps2_kb/_0284_ ) );
BUF_X2 \u0_ps2_kb/_0534_ ( .A(\u0_ps2_kb/_0284_ ), .Z(\u0_ps2_kb/_0285_ ) );
AND2_X1 \u0_ps2_kb/_0535_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0286_ ) );
NAND2_X1 \u0_ps2_kb/_0536_ ( .A1(\u0_ps2_kb/_0282_ ), .A2(\u0_ps2_kb/_0286_ ), .ZN(\u0_ps2_kb/_0287_ ) );
MUX2_X1 \u0_ps2_kb/_0537_ ( .A(\u0_ps2_kb/_0441_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0287_ ), .Z(\u0_ps2_kb/_0102_ ) );
INV_X1 \u0_ps2_kb/_0538_ ( .A(\u0_ps2_kb/_0441_ ), .ZN(\u0_ps2_kb/_0288_ ) );
XOR2_X2 \u0_ps2_kb/_0539_ ( .A(\u0_ps2_kb/_0200_ ), .B(\u0_ps2_kb/_0199_ ), .Z(\u0_ps2_kb/_0289_ ) );
XNOR2_X2 \u0_ps2_kb/_0540_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0193_ ), .ZN(\u0_ps2_kb/_0290_ ) );
XNOR2_X2 \u0_ps2_kb/_0541_ ( .A(\u0_ps2_kb/_0289_ ), .B(\u0_ps2_kb/_0290_ ), .ZN(\u0_ps2_kb/_0291_ ) );
XNOR2_X1 \u0_ps2_kb/_0542_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0197_ ), .ZN(\u0_ps2_kb/_0292_ ) );
XNOR2_X2 \u0_ps2_kb/_0543_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0195_ ), .ZN(\u0_ps2_kb/_0293_ ) );
XNOR2_X1 \u0_ps2_kb/_0544_ ( .A(\u0_ps2_kb/_0292_ ), .B(\u0_ps2_kb/_0293_ ), .ZN(\u0_ps2_kb/_0294_ ) );
XNOR2_X2 \u0_ps2_kb/_0545_ ( .A(\u0_ps2_kb/_0291_ ), .B(\u0_ps2_kb/_0294_ ), .ZN(\u0_ps2_kb/_0295_ ) );
AOI211_X2 \u0_ps2_kb/_0546_ ( .A(\u0_ps2_kb/_0288_ ), .B(\u0_ps2_kb/_0192_ ), .C1(\u0_ps2_kb/_0295_ ), .C2(\u0_ps2_kb/_0201_ ), .ZN(\u0_ps2_kb/_0296_ ) );
OR2_X1 \u0_ps2_kb/_0547_ ( .A1(\u0_ps2_kb/_0295_ ), .A2(\u0_ps2_kb/_0201_ ), .ZN(\u0_ps2_kb/_0297_ ) );
AND2_X2 \u0_ps2_kb/_0548_ ( .A1(\u0_ps2_kb/_0296_ ), .A2(\u0_ps2_kb/_0297_ ), .ZN(\u0_ps2_kb/_0298_ ) );
NOR2_X1 \u0_ps2_kb/_0549_ ( .A1(\u0_ps2_kb/_0281_ ), .A2(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0299_ ) );
AND2_X1 \u0_ps2_kb/_0550_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0299_ ), .ZN(\u0_ps2_kb/_0300_ ) );
AND2_X1 \u0_ps2_kb/_0551_ ( .A1(\u0_ps2_kb/_0300_ ), .A2(\u0_ps2_kb/_0284_ ), .ZN(\u0_ps2_kb/_0301_ ) );
AND2_X4 \u0_ps2_kb/_0552_ ( .A1(\u0_ps2_kb/_0298_ ), .A2(\u0_ps2_kb/_0301_ ), .ZN(\u0_ps2_kb/_0302_ ) );
AND2_X4 \u0_ps2_kb/_0553_ ( .A1(\u0_ps2_kb/_0302_ ), .A2(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0303_ ) );
AND3_X1 \u0_ps2_kb/_0554_ ( .A1(\u0_ps2_kb/_0448_ ), .A2(\u0_ps2_kb/_0447_ ), .A3(\u0_ps2_kb/_0446_ ), .ZN(\u0_ps2_kb/_0304_ ) );
NAND2_X2 \u0_ps2_kb/_0555_ ( .A1(\u0_ps2_kb/_0303_ ), .A2(\u0_ps2_kb/_0304_ ), .ZN(\u0_ps2_kb/_0305_ ) );
MUX2_X1 \u0_ps2_kb/_0556_ ( .A(\u0_ps2_kb/_0193_ ), .B(\u0_ps2_kb/_0271_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0174_ ) );
MUX2_X1 \u0_ps2_kb/_0557_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0272_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0175_ ) );
MUX2_X1 \u0_ps2_kb/_0558_ ( .A(\u0_ps2_kb/_0195_ ), .B(\u0_ps2_kb/_0273_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0176_ ) );
MUX2_X1 \u0_ps2_kb/_0559_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0274_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0177_ ) );
MUX2_X1 \u0_ps2_kb/_0560_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0275_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0178_ ) );
MUX2_X1 \u0_ps2_kb/_0561_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0276_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0179_ ) );
MUX2_X1 \u0_ps2_kb/_0562_ ( .A(\u0_ps2_kb/_0199_ ), .B(\u0_ps2_kb/_0277_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0180_ ) );
MUX2_X1 \u0_ps2_kb/_0563_ ( .A(\u0_ps2_kb/_0200_ ), .B(\u0_ps2_kb/_0278_ ), .S(\u0_ps2_kb/_0305_ ), .Z(\u0_ps2_kb/_0181_ ) );
INV_X1 \u0_ps2_kb/_0564_ ( .A(\u0_ps2_kb/_0446_ ), .ZN(\u0_ps2_kb/_0306_ ) );
AND3_X1 \u0_ps2_kb/_0565_ ( .A1(\u0_ps2_kb/_0306_ ), .A2(\u0_ps2_kb/_0448_ ), .A3(\u0_ps2_kb/_0447_ ), .ZN(\u0_ps2_kb/_0307_ ) );
NAND2_X2 \u0_ps2_kb/_0566_ ( .A1(\u0_ps2_kb/_0303_ ), .A2(\u0_ps2_kb/_0307_ ), .ZN(\u0_ps2_kb/_0308_ ) );
MUX2_X1 \u0_ps2_kb/_0567_ ( .A(\u0_ps2_kb/_0193_ ), .B(\u0_ps2_kb/_0263_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0166_ ) );
MUX2_X1 \u0_ps2_kb/_0568_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0264_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0167_ ) );
MUX2_X1 \u0_ps2_kb/_0569_ ( .A(\u0_ps2_kb/_0195_ ), .B(\u0_ps2_kb/_0265_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0168_ ) );
MUX2_X1 \u0_ps2_kb/_0570_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0266_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0169_ ) );
MUX2_X1 \u0_ps2_kb/_0571_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0267_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0170_ ) );
MUX2_X1 \u0_ps2_kb/_0572_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0268_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0171_ ) );
MUX2_X1 \u0_ps2_kb/_0573_ ( .A(\u0_ps2_kb/_0199_ ), .B(\u0_ps2_kb/_0269_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0172_ ) );
MUX2_X1 \u0_ps2_kb/_0574_ ( .A(\u0_ps2_kb/_0200_ ), .B(\u0_ps2_kb/_0270_ ), .S(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0173_ ) );
AND3_X1 \u0_ps2_kb/_0575_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0299_ ), .A3(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0309_ ) );
NOR2_X1 \u0_ps2_kb/_0576_ ( .A1(\u0_ps2_kb/_0203_ ), .A2(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0310_ ) );
NAND2_X1 \u0_ps2_kb/_0577_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0310_ ), .ZN(\u0_ps2_kb/_0311_ ) );
MUX2_X1 \u0_ps2_kb/_0578_ ( .A(\u0_ps2_kb/_0441_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0311_ ), .Z(\u0_ps2_kb/_0104_ ) );
AND2_X1 \u0_ps2_kb/_0579_ ( .A1(\u0_ps2_kb/_0203_ ), .A2(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0312_ ) );
AND2_X1 \u0_ps2_kb/_0580_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0312_ ), .ZN(\u0_ps2_kb/_0313_ ) );
INV_X1 \u0_ps2_kb/_0581_ ( .A(\u0_ps2_kb/_0313_ ), .ZN(\u0_ps2_kb/_0314_ ) );
NAND3_X1 \u0_ps2_kb/_0582_ ( .A1(\u0_ps2_kb/_0281_ ), .A2(\u0_ps2_kb/_0202_ ), .A3(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0315_ ) );
NOR2_X1 \u0_ps2_kb/_0583_ ( .A1(\u0_ps2_kb/_0314_ ), .A2(\u0_ps2_kb/_0315_ ), .ZN(\u0_ps2_kb/_0316_ ) );
MUX2_X1 \u0_ps2_kb/_0584_ ( .A(\u0_ps2_kb/_0199_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0316_ ), .Z(\u0_ps2_kb/_0103_ ) );
INV_X1 \u0_ps2_kb/_0585_ ( .A(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0317_ ) );
NOR2_X1 \u0_ps2_kb/_0586_ ( .A1(\u0_ps2_kb/_0317_ ), .A2(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0318_ ) );
NAND2_X1 \u0_ps2_kb/_0587_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0318_ ), .ZN(\u0_ps2_kb/_0319_ ) );
MUX2_X1 \u0_ps2_kb/_0588_ ( .A(\u0_ps2_kb/_0441_ ), .B(\u0_ps2_kb/_0201_ ), .S(\u0_ps2_kb/_0319_ ), .Z(\u0_ps2_kb/_0105_ ) );
INV_X1 \u0_ps2_kb/_0589_ ( .A(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0320_ ) );
NOR2_X1 \u0_ps2_kb/_0590_ ( .A1(\u0_ps2_kb/_0320_ ), .A2(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0321_ ) );
NAND2_X1 \u0_ps2_kb/_0591_ ( .A1(\u0_ps2_kb/_0321_ ), .A2(\u0_ps2_kb/_0281_ ), .ZN(\u0_ps2_kb/_0322_ ) );
NOR2_X1 \u0_ps2_kb/_0592_ ( .A1(\u0_ps2_kb/_0314_ ), .A2(\u0_ps2_kb/_0322_ ), .ZN(\u0_ps2_kb/_0323_ ) );
MUX2_X1 \u0_ps2_kb/_0593_ ( .A(\u0_ps2_kb/_0195_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0323_ ), .Z(\u0_ps2_kb/_0099_ ) );
NAND2_X1 \u0_ps2_kb/_0594_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0310_ ), .ZN(\u0_ps2_kb/_0324_ ) );
NOR2_X1 \u0_ps2_kb/_0595_ ( .A1(\u0_ps2_kb/_0324_ ), .A2(\u0_ps2_kb/_0315_ ), .ZN(\u0_ps2_kb/_0325_ ) );
MUX2_X1 \u0_ps2_kb/_0596_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0325_ ), .Z(\u0_ps2_kb/_0100_ ) );
NAND2_X1 \u0_ps2_kb/_0597_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0318_ ), .ZN(\u0_ps2_kb/_0326_ ) );
NOR2_X1 \u0_ps2_kb/_0598_ ( .A1(\u0_ps2_kb/_0326_ ), .A2(\u0_ps2_kb/_0315_ ), .ZN(\u0_ps2_kb/_0327_ ) );
MUX2_X1 \u0_ps2_kb/_0599_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0327_ ), .Z(\u0_ps2_kb/_0101_ ) );
AND2_X4 \u0_ps2_kb/_0600_ ( .A1(\u0_ps2_kb/_0303_ ), .A2(\u0_ps2_kb/_0306_ ), .ZN(\u0_ps2_kb/_0328_ ) );
INV_X1 \u0_ps2_kb/_0601_ ( .A(\u0_ps2_kb/_0448_ ), .ZN(\u0_ps2_kb/_0329_ ) );
NOR2_X1 \u0_ps2_kb/_0602_ ( .A1(\u0_ps2_kb/_0329_ ), .A2(\u0_ps2_kb/_0447_ ), .ZN(\u0_ps2_kb/_0330_ ) );
NAND2_X4 \u0_ps2_kb/_0603_ ( .A1(\u0_ps2_kb/_0328_ ), .A2(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0331_ ) );
MUX2_X1 \u0_ps2_kb/_0604_ ( .A(\u0_ps2_kb/_0193_ ), .B(\u0_ps2_kb/_0247_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0150_ ) );
MUX2_X1 \u0_ps2_kb/_0605_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0248_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0151_ ) );
MUX2_X1 \u0_ps2_kb/_0606_ ( .A(\u0_ps2_kb/_0195_ ), .B(\u0_ps2_kb/_0249_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0152_ ) );
MUX2_X1 \u0_ps2_kb/_0607_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0250_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0153_ ) );
MUX2_X1 \u0_ps2_kb/_0608_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0251_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0154_ ) );
MUX2_X1 \u0_ps2_kb/_0609_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0252_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0155_ ) );
MUX2_X1 \u0_ps2_kb/_0610_ ( .A(\u0_ps2_kb/_0199_ ), .B(\u0_ps2_kb/_0253_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0156_ ) );
MUX2_X1 \u0_ps2_kb/_0611_ ( .A(\u0_ps2_kb/_0200_ ), .B(\u0_ps2_kb/_0254_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0157_ ) );
MUX2_X1 \u0_ps2_kb/_0612_ ( .A(\u0_ps2_kb/_0231_ ), .B(\u0_ps2_kb/_0239_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0332_ ) );
MUX2_X1 \u0_ps2_kb/_0613_ ( .A(\u0_ps2_kb/_0215_ ), .B(\u0_ps2_kb/_0223_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0333_ ) );
INV_X1 \u0_ps2_kb/_0614_ ( .A(\u0_ps2_kb/_0443_ ), .ZN(\u0_ps2_kb/_0334_ ) );
MUX2_X1 \u0_ps2_kb/_0615_ ( .A(\u0_ps2_kb/_0332_ ), .B(\u0_ps2_kb/_0333_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0335_ ) );
MUX2_X1 \u0_ps2_kb/_0616_ ( .A(\u0_ps2_kb/_0247_ ), .B(\u0_ps2_kb/_0263_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0336_ ) );
MUX2_X1 \u0_ps2_kb/_0617_ ( .A(\u0_ps2_kb/_0255_ ), .B(\u0_ps2_kb/_0271_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0337_ ) );
MUX2_X1 \u0_ps2_kb/_0618_ ( .A(\u0_ps2_kb/_0336_ ), .B(\u0_ps2_kb/_0337_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0338_ ) );
MUX2_X1 \u0_ps2_kb/_0619_ ( .A(\u0_ps2_kb/_0335_ ), .B(\u0_ps2_kb/_0338_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0207_ ) );
MUX2_X1 \u0_ps2_kb/_0620_ ( .A(\u0_ps2_kb/_0232_ ), .B(\u0_ps2_kb/_0240_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0339_ ) );
MUX2_X1 \u0_ps2_kb/_0621_ ( .A(\u0_ps2_kb/_0216_ ), .B(\u0_ps2_kb/_0224_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0340_ ) );
MUX2_X1 \u0_ps2_kb/_0622_ ( .A(\u0_ps2_kb/_0339_ ), .B(\u0_ps2_kb/_0340_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0341_ ) );
MUX2_X1 \u0_ps2_kb/_0623_ ( .A(\u0_ps2_kb/_0248_ ), .B(\u0_ps2_kb/_0264_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0342_ ) );
MUX2_X1 \u0_ps2_kb/_0624_ ( .A(\u0_ps2_kb/_0256_ ), .B(\u0_ps2_kb/_0272_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0343_ ) );
MUX2_X1 \u0_ps2_kb/_0625_ ( .A(\u0_ps2_kb/_0342_ ), .B(\u0_ps2_kb/_0343_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0344_ ) );
MUX2_X1 \u0_ps2_kb/_0626_ ( .A(\u0_ps2_kb/_0341_ ), .B(\u0_ps2_kb/_0344_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0208_ ) );
MUX2_X1 \u0_ps2_kb/_0627_ ( .A(\u0_ps2_kb/_0233_ ), .B(\u0_ps2_kb/_0241_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0345_ ) );
MUX2_X1 \u0_ps2_kb/_0628_ ( .A(\u0_ps2_kb/_0217_ ), .B(\u0_ps2_kb/_0225_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0346_ ) );
MUX2_X1 \u0_ps2_kb/_0629_ ( .A(\u0_ps2_kb/_0345_ ), .B(\u0_ps2_kb/_0346_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0347_ ) );
MUX2_X1 \u0_ps2_kb/_0630_ ( .A(\u0_ps2_kb/_0249_ ), .B(\u0_ps2_kb/_0265_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0348_ ) );
MUX2_X1 \u0_ps2_kb/_0631_ ( .A(\u0_ps2_kb/_0257_ ), .B(\u0_ps2_kb/_0273_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0349_ ) );
MUX2_X1 \u0_ps2_kb/_0632_ ( .A(\u0_ps2_kb/_0348_ ), .B(\u0_ps2_kb/_0349_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0350_ ) );
MUX2_X1 \u0_ps2_kb/_0633_ ( .A(\u0_ps2_kb/_0347_ ), .B(\u0_ps2_kb/_0350_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0209_ ) );
MUX2_X1 \u0_ps2_kb/_0634_ ( .A(\u0_ps2_kb/_0234_ ), .B(\u0_ps2_kb/_0242_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0351_ ) );
MUX2_X1 \u0_ps2_kb/_0635_ ( .A(\u0_ps2_kb/_0218_ ), .B(\u0_ps2_kb/_0226_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0352_ ) );
MUX2_X1 \u0_ps2_kb/_0636_ ( .A(\u0_ps2_kb/_0351_ ), .B(\u0_ps2_kb/_0352_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0353_ ) );
MUX2_X1 \u0_ps2_kb/_0637_ ( .A(\u0_ps2_kb/_0250_ ), .B(\u0_ps2_kb/_0266_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0354_ ) );
MUX2_X1 \u0_ps2_kb/_0638_ ( .A(\u0_ps2_kb/_0258_ ), .B(\u0_ps2_kb/_0274_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0355_ ) );
MUX2_X1 \u0_ps2_kb/_0639_ ( .A(\u0_ps2_kb/_0354_ ), .B(\u0_ps2_kb/_0355_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0356_ ) );
MUX2_X1 \u0_ps2_kb/_0640_ ( .A(\u0_ps2_kb/_0353_ ), .B(\u0_ps2_kb/_0356_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0210_ ) );
MUX2_X1 \u0_ps2_kb/_0641_ ( .A(\u0_ps2_kb/_0235_ ), .B(\u0_ps2_kb/_0243_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0357_ ) );
MUX2_X1 \u0_ps2_kb/_0642_ ( .A(\u0_ps2_kb/_0219_ ), .B(\u0_ps2_kb/_0227_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0358_ ) );
MUX2_X1 \u0_ps2_kb/_0643_ ( .A(\u0_ps2_kb/_0357_ ), .B(\u0_ps2_kb/_0358_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0359_ ) );
MUX2_X1 \u0_ps2_kb/_0644_ ( .A(\u0_ps2_kb/_0251_ ), .B(\u0_ps2_kb/_0267_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0360_ ) );
MUX2_X1 \u0_ps2_kb/_0645_ ( .A(\u0_ps2_kb/_0259_ ), .B(\u0_ps2_kb/_0275_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0361_ ) );
MUX2_X1 \u0_ps2_kb/_0646_ ( .A(\u0_ps2_kb/_0360_ ), .B(\u0_ps2_kb/_0361_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0362_ ) );
MUX2_X1 \u0_ps2_kb/_0647_ ( .A(\u0_ps2_kb/_0359_ ), .B(\u0_ps2_kb/_0362_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0211_ ) );
MUX2_X1 \u0_ps2_kb/_0648_ ( .A(\u0_ps2_kb/_0236_ ), .B(\u0_ps2_kb/_0244_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0363_ ) );
MUX2_X1 \u0_ps2_kb/_0649_ ( .A(\u0_ps2_kb/_0220_ ), .B(\u0_ps2_kb/_0228_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0364_ ) );
MUX2_X1 \u0_ps2_kb/_0650_ ( .A(\u0_ps2_kb/_0363_ ), .B(\u0_ps2_kb/_0364_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0365_ ) );
MUX2_X1 \u0_ps2_kb/_0651_ ( .A(\u0_ps2_kb/_0252_ ), .B(\u0_ps2_kb/_0268_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0366_ ) );
MUX2_X1 \u0_ps2_kb/_0652_ ( .A(\u0_ps2_kb/_0260_ ), .B(\u0_ps2_kb/_0276_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0367_ ) );
MUX2_X1 \u0_ps2_kb/_0653_ ( .A(\u0_ps2_kb/_0366_ ), .B(\u0_ps2_kb/_0367_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0368_ ) );
MUX2_X1 \u0_ps2_kb/_0654_ ( .A(\u0_ps2_kb/_0365_ ), .B(\u0_ps2_kb/_0368_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0212_ ) );
MUX2_X1 \u0_ps2_kb/_0655_ ( .A(\u0_ps2_kb/_0221_ ), .B(\u0_ps2_kb/_0237_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0369_ ) );
MUX2_X1 \u0_ps2_kb/_0656_ ( .A(\u0_ps2_kb/_0229_ ), .B(\u0_ps2_kb/_0245_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0370_ ) );
MUX2_X1 \u0_ps2_kb/_0657_ ( .A(\u0_ps2_kb/_0369_ ), .B(\u0_ps2_kb/_0370_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0371_ ) );
MUX2_X1 \u0_ps2_kb/_0658_ ( .A(\u0_ps2_kb/_0253_ ), .B(\u0_ps2_kb/_0269_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0372_ ) );
MUX2_X1 \u0_ps2_kb/_0659_ ( .A(\u0_ps2_kb/_0261_ ), .B(\u0_ps2_kb/_0277_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0373_ ) );
MUX2_X1 \u0_ps2_kb/_0660_ ( .A(\u0_ps2_kb/_0372_ ), .B(\u0_ps2_kb/_0373_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0374_ ) );
MUX2_X1 \u0_ps2_kb/_0661_ ( .A(\u0_ps2_kb/_0371_ ), .B(\u0_ps2_kb/_0374_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0213_ ) );
MUX2_X1 \u0_ps2_kb/_0662_ ( .A(\u0_ps2_kb/_0238_ ), .B(\u0_ps2_kb/_0246_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0375_ ) );
MUX2_X1 \u0_ps2_kb/_0663_ ( .A(\u0_ps2_kb/_0222_ ), .B(\u0_ps2_kb/_0230_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0376_ ) );
MUX2_X1 \u0_ps2_kb/_0664_ ( .A(\u0_ps2_kb/_0375_ ), .B(\u0_ps2_kb/_0376_ ), .S(\u0_ps2_kb/_0334_ ), .Z(\u0_ps2_kb/_0377_ ) );
MUX2_X1 \u0_ps2_kb/_0665_ ( .A(\u0_ps2_kb/_0254_ ), .B(\u0_ps2_kb/_0270_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0378_ ) );
MUX2_X1 \u0_ps2_kb/_0666_ ( .A(\u0_ps2_kb/_0262_ ), .B(\u0_ps2_kb/_0278_ ), .S(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0379_ ) );
MUX2_X1 \u0_ps2_kb/_0667_ ( .A(\u0_ps2_kb/_0378_ ), .B(\u0_ps2_kb/_0379_ ), .S(\u0_ps2_kb/_0442_ ), .Z(\u0_ps2_kb/_0380_ ) );
MUX2_X1 \u0_ps2_kb/_0668_ ( .A(\u0_ps2_kb/_0377_ ), .B(\u0_ps2_kb/_0380_ ), .S(\u0_ps2_kb/_0444_ ), .Z(\u0_ps2_kb/_0214_ ) );
INV_X1 \u0_ps2_kb/_0669_ ( .A(\u0_ps2_kb/_0184_ ), .ZN(\u0_ps2_kb/_0381_ ) );
AND3_X2 \u0_ps2_kb/_0670_ ( .A1(\u0_ps2_kb/_0298_ ), .A2(\u0_ps2_kb/_0381_ ), .A3(\u0_ps2_kb/_0301_ ), .ZN(\u0_ps2_kb/_0382_ ) );
NAND2_X2 \u0_ps2_kb/_0671_ ( .A1(\u0_ps2_kb/_0382_ ), .A2(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0383_ ) );
NAND2_X1 \u0_ps2_kb/_0672_ ( .A1(\u0_ps2_kb/_0329_ ), .A2(\u0_ps2_kb/_0447_ ), .ZN(\u0_ps2_kb/_0384_ ) );
NOR2_X4 \u0_ps2_kb/_0673_ ( .A1(\u0_ps2_kb/_0383_ ), .A2(\u0_ps2_kb/_0384_ ), .ZN(\u0_ps2_kb/_0385_ ) );
MUX2_X1 \u0_ps2_kb/_0674_ ( .A(\u0_ps2_kb/_0239_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0142_ ) );
MUX2_X1 \u0_ps2_kb/_0675_ ( .A(\u0_ps2_kb/_0240_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0143_ ) );
MUX2_X1 \u0_ps2_kb/_0676_ ( .A(\u0_ps2_kb/_0241_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0144_ ) );
MUX2_X1 \u0_ps2_kb/_0677_ ( .A(\u0_ps2_kb/_0242_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0145_ ) );
MUX2_X1 \u0_ps2_kb/_0678_ ( .A(\u0_ps2_kb/_0243_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0146_ ) );
MUX2_X1 \u0_ps2_kb/_0679_ ( .A(\u0_ps2_kb/_0244_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0147_ ) );
MUX2_X1 \u0_ps2_kb/_0680_ ( .A(\u0_ps2_kb/_0245_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0148_ ) );
MUX2_X1 \u0_ps2_kb/_0681_ ( .A(\u0_ps2_kb/_0246_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0385_ ), .Z(\u0_ps2_kb/_0149_ ) );
INV_X4 \u0_ps2_kb/_0682_ ( .A(\u0_ps2_kb/_0328_ ), .ZN(\u0_ps2_kb/_0386_ ) );
NOR2_X4 \u0_ps2_kb/_0683_ ( .A1(\u0_ps2_kb/_0386_ ), .A2(\u0_ps2_kb/_0384_ ), .ZN(\u0_ps2_kb/_0387_ ) );
MUX2_X1 \u0_ps2_kb/_0684_ ( .A(\u0_ps2_kb/_0231_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0134_ ) );
MUX2_X1 \u0_ps2_kb/_0685_ ( .A(\u0_ps2_kb/_0232_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0135_ ) );
MUX2_X1 \u0_ps2_kb/_0686_ ( .A(\u0_ps2_kb/_0233_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0136_ ) );
MUX2_X1 \u0_ps2_kb/_0687_ ( .A(\u0_ps2_kb/_0234_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0137_ ) );
MUX2_X1 \u0_ps2_kb/_0688_ ( .A(\u0_ps2_kb/_0235_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0138_ ) );
MUX2_X1 \u0_ps2_kb/_0689_ ( .A(\u0_ps2_kb/_0236_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0139_ ) );
MUX2_X1 \u0_ps2_kb/_0690_ ( .A(\u0_ps2_kb/_0237_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0140_ ) );
MUX2_X1 \u0_ps2_kb/_0691_ ( .A(\u0_ps2_kb/_0238_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0387_ ), .Z(\u0_ps2_kb/_0141_ ) );
OR2_X1 \u0_ps2_kb/_0692_ ( .A1(\u0_ps2_kb/_0448_ ), .A2(\u0_ps2_kb/_0447_ ), .ZN(\u0_ps2_kb/_0388_ ) );
NOR2_X4 \u0_ps2_kb/_0693_ ( .A1(\u0_ps2_kb/_0383_ ), .A2(\u0_ps2_kb/_0388_ ), .ZN(\u0_ps2_kb/_0389_ ) );
MUX2_X1 \u0_ps2_kb/_0694_ ( .A(\u0_ps2_kb/_0223_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0126_ ) );
MUX2_X1 \u0_ps2_kb/_0695_ ( .A(\u0_ps2_kb/_0224_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0127_ ) );
MUX2_X1 \u0_ps2_kb/_0696_ ( .A(\u0_ps2_kb/_0225_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0128_ ) );
MUX2_X1 \u0_ps2_kb/_0697_ ( .A(\u0_ps2_kb/_0226_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0129_ ) );
MUX2_X1 \u0_ps2_kb/_0698_ ( .A(\u0_ps2_kb/_0227_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0130_ ) );
MUX2_X1 \u0_ps2_kb/_0699_ ( .A(\u0_ps2_kb/_0228_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0131_ ) );
MUX2_X1 \u0_ps2_kb/_0700_ ( .A(\u0_ps2_kb/_0229_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0132_ ) );
MUX2_X1 \u0_ps2_kb/_0701_ ( .A(\u0_ps2_kb/_0230_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0389_ ), .Z(\u0_ps2_kb/_0133_ ) );
NOR2_X4 \u0_ps2_kb/_0702_ ( .A1(\u0_ps2_kb/_0386_ ), .A2(\u0_ps2_kb/_0388_ ), .ZN(\u0_ps2_kb/_0390_ ) );
MUX2_X1 \u0_ps2_kb/_0703_ ( .A(\u0_ps2_kb/_0215_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0118_ ) );
MUX2_X1 \u0_ps2_kb/_0704_ ( .A(\u0_ps2_kb/_0216_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0119_ ) );
MUX2_X1 \u0_ps2_kb/_0705_ ( .A(\u0_ps2_kb/_0217_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0120_ ) );
MUX2_X1 \u0_ps2_kb/_0706_ ( .A(\u0_ps2_kb/_0218_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0121_ ) );
MUX2_X1 \u0_ps2_kb/_0707_ ( .A(\u0_ps2_kb/_0219_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0122_ ) );
MUX2_X1 \u0_ps2_kb/_0708_ ( .A(\u0_ps2_kb/_0220_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0123_ ) );
MUX2_X1 \u0_ps2_kb/_0709_ ( .A(\u0_ps2_kb/_0221_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0124_ ) );
MUX2_X1 \u0_ps2_kb/_0710_ ( .A(\u0_ps2_kb/_0222_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0390_ ), .Z(\u0_ps2_kb/_0125_ ) );
NAND2_X1 \u0_ps2_kb/_0711_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0285_ ), .ZN(\u0_ps2_kb/_0391_ ) );
NOR2_X1 \u0_ps2_kb/_0712_ ( .A1(\u0_ps2_kb/_0391_ ), .A2(\u0_ps2_kb/_0322_ ), .ZN(\u0_ps2_kb/_0392_ ) );
MUX2_X1 \u0_ps2_kb/_0713_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0392_ ), .Z(\u0_ps2_kb/_0098_ ) );
NOR2_X1 \u0_ps2_kb/_0714_ ( .A1(\u0_ps2_kb/_0326_ ), .A2(\u0_ps2_kb/_0322_ ), .ZN(\u0_ps2_kb/_0393_ ) );
MUX2_X1 \u0_ps2_kb/_0715_ ( .A(\u0_ps2_kb/_0193_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0393_ ), .Z(\u0_ps2_kb/_0097_ ) );
NOR2_X1 \u0_ps2_kb/_0716_ ( .A1(\u0_ps2_kb/_0324_ ), .A2(\u0_ps2_kb/_0322_ ), .ZN(\u0_ps2_kb/_0394_ ) );
MUX2_X1 \u0_ps2_kb/_0717_ ( .A(\u0_ps2_kb/_0192_ ), .B(\u0_ps2_kb/_0441_ ), .S(\u0_ps2_kb/_0394_ ), .Z(\u0_ps2_kb/_0096_ ) );
BUF_X4 \u0_ps2_kb/_0718_ ( .A(\u0_ps2_kb/_0320_ ), .Z(\u0_ps2_kb/_0395_ ) );
XNOR2_X1 \u0_ps2_kb/_0719_ ( .A(\u0_ps2_kb/_0285_ ), .B(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0396_ ) );
NOR3_X1 \u0_ps2_kb/_0720_ ( .A1(\u0_ps2_kb/_0301_ ), .A2(\u0_ps2_kb/_0395_ ), .A3(\u0_ps2_kb/_0396_ ), .ZN(\u0_ps2_kb/_0106_ ) );
NOR3_X1 \u0_ps2_kb/_0721_ ( .A1(\u0_ps2_kb/_0299_ ), .A2(\u0_ps2_kb/_0203_ ), .A3(\u0_ps2_kb/_0279_ ), .ZN(\u0_ps2_kb/_0397_ ) );
INV_X1 \u0_ps2_kb/_0722_ ( .A(\u0_ps2_kb/_0285_ ), .ZN(\u0_ps2_kb/_0398_ ) );
NOR3_X1 \u0_ps2_kb/_0723_ ( .A1(\u0_ps2_kb/_0397_ ), .A2(\u0_ps2_kb/_0398_ ), .A3(\u0_ps2_kb/_0318_ ), .ZN(\u0_ps2_kb/_0399_ ) );
AOI211_X4 \u0_ps2_kb/_0724_ ( .A(\u0_ps2_kb/_0395_ ), .B(\u0_ps2_kb/_0399_ ), .C1(\u0_ps2_kb/_0185_ ), .C2(\u0_ps2_kb/_0398_ ), .ZN(\u0_ps2_kb/_0107_ ) );
XNOR2_X1 \u0_ps2_kb/_0725_ ( .A(\u0_ps2_kb/_0313_ ), .B(\u0_ps2_kb/_0186_ ), .ZN(\u0_ps2_kb/_0400_ ) );
INV_X1 \u0_ps2_kb/_0726_ ( .A(\u0_ps2_kb/_0301_ ), .ZN(\u0_ps2_kb/_0401_ ) );
AND3_X1 \u0_ps2_kb/_0727_ ( .A1(\u0_ps2_kb/_0400_ ), .A2(\u0_ps2_kb/_0202_ ), .A3(\u0_ps2_kb/_0401_ ), .ZN(\u0_ps2_kb/_0108_ ) );
NAND3_X1 \u0_ps2_kb/_0728_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0205_ ), .A3(\u0_ps2_kb/_0312_ ), .ZN(\u0_ps2_kb/_0402_ ) );
OAI211_X2 \u0_ps2_kb/_0729_ ( .A(\u0_ps2_kb/_0401_ ), .B(\u0_ps2_kb/_0202_ ), .C1(\u0_ps2_kb/_0187_ ), .C2(\u0_ps2_kb/_0402_ ), .ZN(\u0_ps2_kb/_0403_ ) );
AOI21_X1 \u0_ps2_kb/_0730_ ( .A(\u0_ps2_kb/_0403_ ), .B1(\u0_ps2_kb/_0187_ ), .B2(\u0_ps2_kb/_0402_ ), .ZN(\u0_ps2_kb/_0109_ ) );
XNOR2_X1 \u0_ps2_kb/_0731_ ( .A(\u0_ps2_kb/_0442_ ), .B(\u0_ps2_kb/_0437_ ), .ZN(\u0_ps2_kb/_0404_ ) );
NAND2_X1 \u0_ps2_kb/_0732_ ( .A1(\u0_ps2_kb/_0404_ ), .A2(\u0_ps2_kb/_0445_ ), .ZN(\u0_ps2_kb/_0405_ ) );
OR2_X1 \u0_ps2_kb/_0733_ ( .A1(\u0_ps2_kb/_0188_ ), .A2(\u0_ps2_kb/_0445_ ), .ZN(\u0_ps2_kb/_0406_ ) );
AOI21_X1 \u0_ps2_kb/_0734_ ( .A(\u0_ps2_kb/_0395_ ), .B1(\u0_ps2_kb/_0405_ ), .B2(\u0_ps2_kb/_0406_ ), .ZN(\u0_ps2_kb/_0111_ ) );
XOR2_X1 \u0_ps2_kb/_0735_ ( .A(\u0_ps2_kb/_0442_ ), .B(\u0_ps2_kb/_0443_ ), .Z(\u0_ps2_kb/_0407_ ) );
INV_X1 \u0_ps2_kb/_0736_ ( .A(\u0_ps2_kb/_0437_ ), .ZN(\u0_ps2_kb/_0408_ ) );
NAND2_X1 \u0_ps2_kb/_0737_ ( .A1(\u0_ps2_kb/_0408_ ), .A2(\u0_ps2_kb/_0445_ ), .ZN(\u0_ps2_kb/_0409_ ) );
NOR2_X1 \u0_ps2_kb/_0738_ ( .A1(\u0_ps2_kb/_0407_ ), .A2(\u0_ps2_kb/_0409_ ), .ZN(\u0_ps2_kb/_0410_ ) );
AOI211_X4 \u0_ps2_kb/_0739_ ( .A(\u0_ps2_kb/_0395_ ), .B(\u0_ps2_kb/_0410_ ), .C1(\u0_ps2_kb/_0183_ ), .C2(\u0_ps2_kb/_0409_ ), .ZN(\u0_ps2_kb/_0112_ ) );
NAND2_X1 \u0_ps2_kb/_0740_ ( .A1(\u0_ps2_kb/_0442_ ), .A2(\u0_ps2_kb/_0443_ ), .ZN(\u0_ps2_kb/_0411_ ) );
XNOR2_X1 \u0_ps2_kb/_0741_ ( .A(\u0_ps2_kb/_0411_ ), .B(\u0_ps2_kb/_0182_ ), .ZN(\u0_ps2_kb/_0412_ ) );
AND3_X1 \u0_ps2_kb/_0742_ ( .A1(\u0_ps2_kb/_0412_ ), .A2(\u0_ps2_kb/_0408_ ), .A3(\u0_ps2_kb/_0445_ ), .ZN(\u0_ps2_kb/_0413_ ) );
AOI211_X4 \u0_ps2_kb/_0743_ ( .A(\u0_ps2_kb/_0395_ ), .B(\u0_ps2_kb/_0413_ ), .C1(\u0_ps2_kb/_0182_ ), .C2(\u0_ps2_kb/_0409_ ), .ZN(\u0_ps2_kb/_0113_ ) );
AOI21_X1 \u0_ps2_kb/_0744_ ( .A(\u0_ps2_kb/_0381_ ), .B1(\u0_ps2_kb/_0298_ ), .B2(\u0_ps2_kb/_0301_ ), .ZN(\u0_ps2_kb/_0414_ ) );
NOR3_X1 \u0_ps2_kb/_0745_ ( .A1(\u0_ps2_kb/_0382_ ), .A2(\u0_ps2_kb/_0414_ ), .A3(\u0_ps2_kb/_0395_ ), .ZN(\u0_ps2_kb/_0115_ ) );
AND2_X1 \u0_ps2_kb/_0746_ ( .A1(\u0_ps2_kb/_0298_ ), .A2(\u0_ps2_kb/_0300_ ), .ZN(\u0_ps2_kb/_0415_ ) );
INV_X1 \u0_ps2_kb/_0747_ ( .A(\u0_ps2_kb/_0415_ ), .ZN(\u0_ps2_kb/_0416_ ) );
XNOR2_X1 \u0_ps2_kb/_0748_ ( .A(\u0_ps2_kb/_0447_ ), .B(\u0_ps2_kb/_0446_ ), .ZN(\u0_ps2_kb/_0417_ ) );
NOR2_X2 \u0_ps2_kb/_0749_ ( .A1(\u0_ps2_kb/_0416_ ), .A2(\u0_ps2_kb/_0417_ ), .ZN(\u0_ps2_kb/_0418_ ) );
OAI21_X1 \u0_ps2_kb/_0750_ ( .A(\u0_ps2_kb/_0285_ ), .B1(\u0_ps2_kb/_0415_ ), .B2(\u0_ps2_kb/_0189_ ), .ZN(\u0_ps2_kb/_0419_ ) );
NOR2_X1 \u0_ps2_kb/_0751_ ( .A1(\u0_ps2_kb/_0418_ ), .A2(\u0_ps2_kb/_0419_ ), .ZN(\u0_ps2_kb/_0420_ ) );
AOI211_X2 \u0_ps2_kb/_0752_ ( .A(\u0_ps2_kb/_0395_ ), .B(\u0_ps2_kb/_0420_ ), .C1(\u0_ps2_kb/_0189_ ), .C2(\u0_ps2_kb/_0398_ ), .ZN(\u0_ps2_kb/_0116_ ) );
NAND2_X1 \u0_ps2_kb/_0753_ ( .A1(\u0_ps2_kb/_0447_ ), .A2(\u0_ps2_kb/_0446_ ), .ZN(\u0_ps2_kb/_0421_ ) );
XNOR2_X1 \u0_ps2_kb/_0754_ ( .A(\u0_ps2_kb/_0421_ ), .B(\u0_ps2_kb/_0190_ ), .ZN(\u0_ps2_kb/_0422_ ) );
AND4_X1 \u0_ps2_kb/_0755_ ( .A1(\u0_ps2_kb/_0297_ ), .A2(\u0_ps2_kb/_0296_ ), .A3(\u0_ps2_kb/_0301_ ), .A4(\u0_ps2_kb/_0422_ ), .ZN(\u0_ps2_kb/_0423_ ) );
INV_X1 \u0_ps2_kb/_0756_ ( .A(\u0_ps2_kb/_0302_ ), .ZN(\u0_ps2_kb/_0424_ ) );
AOI211_X4 \u0_ps2_kb/_0757_ ( .A(\u0_ps2_kb/_0395_ ), .B(\u0_ps2_kb/_0423_ ), .C1(\u0_ps2_kb/_0424_ ), .C2(\u0_ps2_kb/_0190_ ), .ZN(\u0_ps2_kb/_0117_ ) );
AND3_X1 \u0_ps2_kb/_0758_ ( .A1(\u0_ps2_kb/_0415_ ), .A2(\u0_ps2_kb/_0381_ ), .A3(\u0_ps2_kb/_0286_ ), .ZN(\u0_ps2_kb/_0425_ ) );
NAND2_X2 \u0_ps2_kb/_0759_ ( .A1(\u0_ps2_kb/_0425_ ), .A2(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0426_ ) );
MUX2_X1 \u0_ps2_kb/_0760_ ( .A(\u0_ps2_kb/_0193_ ), .B(\u0_ps2_kb/_0255_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0158_ ) );
MUX2_X1 \u0_ps2_kb/_0761_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0256_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0159_ ) );
MUX2_X1 \u0_ps2_kb/_0762_ ( .A(\u0_ps2_kb/_0195_ ), .B(\u0_ps2_kb/_0257_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0160_ ) );
MUX2_X1 \u0_ps2_kb/_0763_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0258_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0161_ ) );
MUX2_X1 \u0_ps2_kb/_0764_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0259_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0162_ ) );
MUX2_X1 \u0_ps2_kb/_0765_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0260_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0163_ ) );
MUX2_X1 \u0_ps2_kb/_0766_ ( .A(\u0_ps2_kb/_0199_ ), .B(\u0_ps2_kb/_0261_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0164_ ) );
MUX2_X1 \u0_ps2_kb/_0767_ ( .A(\u0_ps2_kb/_0200_ ), .B(\u0_ps2_kb/_0262_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0165_ ) );
XNOR2_X1 \u0_ps2_kb/_0768_ ( .A(\u0_ps2_kb/_0407_ ), .B(\u0_ps2_kb/_0189_ ), .ZN(\u0_ps2_kb/_0427_ ) );
XNOR2_X1 \u0_ps2_kb/_0769_ ( .A(\u0_ps2_kb/_0446_ ), .B(\u0_ps2_kb/_0442_ ), .ZN(\u0_ps2_kb/_0428_ ) );
OR3_X1 \u0_ps2_kb/_0770_ ( .A1(\u0_ps2_kb/_0427_ ), .A2(\u0_ps2_kb/_0437_ ), .A3(\u0_ps2_kb/_0428_ ), .ZN(\u0_ps2_kb/_0429_ ) );
XOR2_X1 \u0_ps2_kb/_0771_ ( .A(\u0_ps2_kb/_0412_ ), .B(\u0_ps2_kb/_0190_ ), .Z(\u0_ps2_kb/_0430_ ) );
OAI211_X2 \u0_ps2_kb/_0772_ ( .A(\u0_ps2_kb/_0202_ ), .B(\u0_ps2_kb/_0445_ ), .C1(\u0_ps2_kb/_0429_ ), .C2(\u0_ps2_kb/_0430_ ), .ZN(\u0_ps2_kb/_0431_ ) );
OAI21_X1 \u0_ps2_kb/_0773_ ( .A(\u0_ps2_kb/_0431_ ), .B1(\u0_ps2_kb/_0424_ ), .B2(\u0_ps2_kb/_0395_ ), .ZN(\u0_ps2_kb/_0114_ ) );
XOR2_X1 \u0_ps2_kb/_0774_ ( .A(\u0_ps2_kb/_0422_ ), .B(\u0_ps2_kb/_0182_ ), .Z(\u0_ps2_kb/_0432_ ) );
XOR2_X1 \u0_ps2_kb/_0775_ ( .A(\u0_ps2_kb/_0417_ ), .B(\u0_ps2_kb/_0183_ ), .Z(\u0_ps2_kb/_0433_ ) );
NOR3_X1 \u0_ps2_kb/_0776_ ( .A1(\u0_ps2_kb/_0432_ ), .A2(\u0_ps2_kb/_0428_ ), .A3(\u0_ps2_kb/_0433_ ), .ZN(\u0_ps2_kb/_0434_ ) );
NAND3_X1 \u0_ps2_kb/_0777_ ( .A1(\u0_ps2_kb/_0296_ ), .A2(\u0_ps2_kb/_0297_ ), .A3(\u0_ps2_kb/_0434_ ), .ZN(\u0_ps2_kb/_0435_ ) );
NOR4_X1 \u0_ps2_kb/_0778_ ( .A1(\u0_ps2_kb/_0391_ ), .A2(\u0_ps2_kb/_0205_ ), .A3(\u0_ps2_kb/_0281_ ), .A4(\u0_ps2_kb/_0438_ ), .ZN(\u0_ps2_kb/_0436_ ) );
AOI221_X4 \u0_ps2_kb/_0779_ ( .A(\u0_ps2_kb/_0395_ ), .B1(\u0_ps2_kb/_0191_ ), .B2(\u0_ps2_kb/_0401_ ), .C1(\u0_ps2_kb/_0435_ ), .C2(\u0_ps2_kb/_0436_ ), .ZN(\u0_ps2_kb/_0110_ ) );
BUF_X1 \u0_ps2_kb/_0780_ ( .A(fanout_net_28 ), .Z(\u0_ps2_kb/_0202_ ) );
BUF_X1 \u0_ps2_kb/_0781_ ( .A(\u0_ps2_kb/ps2_clk_sync [1] ), .Z(\u0_ps2_kb/_0439_ ) );
BUF_X1 \u0_ps2_kb/_0782_ ( .A(\u0_ps2_kb/ps2_clk_sync [2] ), .Z(\u0_ps2_kb/_0440_ ) );
BUF_X1 \u0_ps2_kb/_0783_ ( .A(\u0_ps2_kb/count [0] ), .Z(\u0_ps2_kb/_0203_ ) );
BUF_X1 \u0_ps2_kb/_0784_ ( .A(\u0_ps2_kb/count [1] ), .Z(\u0_ps2_kb/_0204_ ) );
BUF_X1 \u0_ps2_kb/_0785_ ( .A(\u0_ps2_kb/count [2] ), .Z(\u0_ps2_kb/_0205_ ) );
BUF_X1 \u0_ps2_kb/_0786_ ( .A(\u0_ps2_kb/count [3] ), .Z(\u0_ps2_kb/_0206_ ) );
BUF_X1 \u0_ps2_kb/_0787_ ( .A(ps2_data ), .Z(\u0_ps2_kb/_0441_ ) );
BUF_X1 \u0_ps2_kb/_0788_ ( .A(\u0_ps2_kb/buffer [6] ), .Z(\u0_ps2_kb/_0198_ ) );
BUF_X1 \u0_ps2_kb/_0789_ ( .A(\u0_ps2_kb/_0102_ ), .Z(\u0_ps2_kb/_0006_ ) );
BUF_X1 \u0_ps2_kb/_0790_ ( .A(\u0_ps2_kb/w_ptr [2] ), .Z(\u0_ps2_kb/_0448_ ) );
BUF_X1 \u0_ps2_kb/_0791_ ( .A(\u0_ps2_kb/w_ptr [1] ), .Z(\u0_ps2_kb/_0447_ ) );
BUF_X1 \u0_ps2_kb/_0792_ ( .A(\u0_ps2_kb/w_ptr [0] ), .Z(\u0_ps2_kb/_0446_ ) );
BUF_X1 \u0_ps2_kb/_0793_ ( .A(\u0_ps2_kb/buffer [0] ), .Z(\u0_ps2_kb/_0192_ ) );
BUF_X1 \u0_ps2_kb/_0794_ ( .A(\u0_ps2_kb/buffer [2] ), .Z(\u0_ps2_kb/_0194_ ) );
BUF_X1 \u0_ps2_kb/_0795_ ( .A(\u0_ps2_kb/buffer [1] ), .Z(\u0_ps2_kb/_0193_ ) );
BUF_X1 \u0_ps2_kb/_0796_ ( .A(\u0_ps2_kb/buffer [4] ), .Z(\u0_ps2_kb/_0196_ ) );
BUF_X1 \u0_ps2_kb/_0797_ ( .A(\u0_ps2_kb/buffer [3] ), .Z(\u0_ps2_kb/_0195_ ) );
BUF_X1 \u0_ps2_kb/_0798_ ( .A(\u0_ps2_kb/buffer [5] ), .Z(\u0_ps2_kb/_0197_ ) );
BUF_X1 \u0_ps2_kb/_0799_ ( .A(\u0_ps2_kb/buffer [8] ), .Z(\u0_ps2_kb/_0200_ ) );
BUF_X1 \u0_ps2_kb/_0800_ ( .A(\u0_ps2_kb/buffer [7] ), .Z(\u0_ps2_kb/_0199_ ) );
BUF_X1 \u0_ps2_kb/_0801_ ( .A(\u0_ps2_kb/buffer [9] ), .Z(\u0_ps2_kb/_0201_ ) );
BUF_X1 \u0_ps2_kb/_0802_ ( .A(\u0_ps2_kb/fifo[7][0] ), .Z(\u0_ps2_kb/_0271_ ) );
BUF_X1 \u0_ps2_kb/_0803_ ( .A(\u0_ps2_kb/_0174_ ), .Z(\u0_ps2_kb/_0078_ ) );
BUF_X1 \u0_ps2_kb/_0804_ ( .A(\u0_ps2_kb/fifo[7][1] ), .Z(\u0_ps2_kb/_0272_ ) );
BUF_X1 \u0_ps2_kb/_0805_ ( .A(\u0_ps2_kb/_0175_ ), .Z(\u0_ps2_kb/_0079_ ) );
BUF_X1 \u0_ps2_kb/_0806_ ( .A(\u0_ps2_kb/fifo[7][2] ), .Z(\u0_ps2_kb/_0273_ ) );
BUF_X1 \u0_ps2_kb/_0807_ ( .A(\u0_ps2_kb/_0176_ ), .Z(\u0_ps2_kb/_0080_ ) );
BUF_X1 \u0_ps2_kb/_0808_ ( .A(\u0_ps2_kb/fifo[7][3] ), .Z(\u0_ps2_kb/_0274_ ) );
BUF_X1 \u0_ps2_kb/_0809_ ( .A(\u0_ps2_kb/_0177_ ), .Z(\u0_ps2_kb/_0081_ ) );
BUF_X1 \u0_ps2_kb/_0810_ ( .A(\u0_ps2_kb/fifo[7][4] ), .Z(\u0_ps2_kb/_0275_ ) );
BUF_X1 \u0_ps2_kb/_0811_ ( .A(\u0_ps2_kb/_0178_ ), .Z(\u0_ps2_kb/_0082_ ) );
BUF_X1 \u0_ps2_kb/_0812_ ( .A(\u0_ps2_kb/fifo[7][5] ), .Z(\u0_ps2_kb/_0276_ ) );
BUF_X1 \u0_ps2_kb/_0813_ ( .A(\u0_ps2_kb/_0179_ ), .Z(\u0_ps2_kb/_0083_ ) );
BUF_X1 \u0_ps2_kb/_0814_ ( .A(\u0_ps2_kb/fifo[7][6] ), .Z(\u0_ps2_kb/_0277_ ) );
BUF_X1 \u0_ps2_kb/_0815_ ( .A(\u0_ps2_kb/_0180_ ), .Z(\u0_ps2_kb/_0084_ ) );
BUF_X1 \u0_ps2_kb/_0816_ ( .A(\u0_ps2_kb/fifo[7][7] ), .Z(\u0_ps2_kb/_0278_ ) );
BUF_X1 \u0_ps2_kb/_0817_ ( .A(\u0_ps2_kb/_0181_ ), .Z(\u0_ps2_kb/_0085_ ) );
BUF_X1 \u0_ps2_kb/_0818_ ( .A(\u0_ps2_kb/fifo[6][0] ), .Z(\u0_ps2_kb/_0263_ ) );
BUF_X1 \u0_ps2_kb/_0819_ ( .A(\u0_ps2_kb/_0166_ ), .Z(\u0_ps2_kb/_0070_ ) );
BUF_X1 \u0_ps2_kb/_0820_ ( .A(\u0_ps2_kb/fifo[6][1] ), .Z(\u0_ps2_kb/_0264_ ) );
BUF_X1 \u0_ps2_kb/_0821_ ( .A(\u0_ps2_kb/_0167_ ), .Z(\u0_ps2_kb/_0071_ ) );
BUF_X1 \u0_ps2_kb/_0822_ ( .A(\u0_ps2_kb/fifo[6][2] ), .Z(\u0_ps2_kb/_0265_ ) );
BUF_X1 \u0_ps2_kb/_0823_ ( .A(\u0_ps2_kb/_0168_ ), .Z(\u0_ps2_kb/_0072_ ) );
BUF_X1 \u0_ps2_kb/_0824_ ( .A(\u0_ps2_kb/fifo[6][3] ), .Z(\u0_ps2_kb/_0266_ ) );
BUF_X1 \u0_ps2_kb/_0825_ ( .A(\u0_ps2_kb/_0169_ ), .Z(\u0_ps2_kb/_0073_ ) );
BUF_X1 \u0_ps2_kb/_0826_ ( .A(\u0_ps2_kb/fifo[6][4] ), .Z(\u0_ps2_kb/_0267_ ) );
BUF_X1 \u0_ps2_kb/_0827_ ( .A(\u0_ps2_kb/_0170_ ), .Z(\u0_ps2_kb/_0074_ ) );
BUF_X1 \u0_ps2_kb/_0828_ ( .A(\u0_ps2_kb/fifo[6][5] ), .Z(\u0_ps2_kb/_0268_ ) );
BUF_X1 \u0_ps2_kb/_0829_ ( .A(\u0_ps2_kb/_0171_ ), .Z(\u0_ps2_kb/_0075_ ) );
BUF_X1 \u0_ps2_kb/_0830_ ( .A(\u0_ps2_kb/fifo[6][6] ), .Z(\u0_ps2_kb/_0269_ ) );
BUF_X1 \u0_ps2_kb/_0831_ ( .A(\u0_ps2_kb/_0172_ ), .Z(\u0_ps2_kb/_0076_ ) );
BUF_X1 \u0_ps2_kb/_0832_ ( .A(\u0_ps2_kb/fifo[6][7] ), .Z(\u0_ps2_kb/_0270_ ) );
BUF_X1 \u0_ps2_kb/_0833_ ( .A(\u0_ps2_kb/_0173_ ), .Z(\u0_ps2_kb/_0077_ ) );
BUF_X1 \u0_ps2_kb/_0834_ ( .A(\u0_ps2_kb/_0104_ ), .Z(\u0_ps2_kb/_0008_ ) );
BUF_X1 \u0_ps2_kb/_0835_ ( .A(\u0_ps2_kb/_0103_ ), .Z(\u0_ps2_kb/_0007_ ) );
BUF_X1 \u0_ps2_kb/_0836_ ( .A(\u0_ps2_kb/_0105_ ), .Z(\u0_ps2_kb/_0009_ ) );
BUF_X1 \u0_ps2_kb/_0837_ ( .A(\u0_ps2_kb/_0099_ ), .Z(\u0_ps2_kb/_0003_ ) );
BUF_X1 \u0_ps2_kb/_0838_ ( .A(\u0_ps2_kb/_0100_ ), .Z(\u0_ps2_kb/_0004_ ) );
BUF_X1 \u0_ps2_kb/_0839_ ( .A(\u0_ps2_kb/_0101_ ), .Z(\u0_ps2_kb/_0005_ ) );
BUF_X1 \u0_ps2_kb/_0840_ ( .A(\u0_ps2_kb/fifo[4][0] ), .Z(\u0_ps2_kb/_0247_ ) );
BUF_X1 \u0_ps2_kb/_0841_ ( .A(\u0_ps2_kb/_0150_ ), .Z(\u0_ps2_kb/_0054_ ) );
BUF_X1 \u0_ps2_kb/_0842_ ( .A(\u0_ps2_kb/fifo[4][1] ), .Z(\u0_ps2_kb/_0248_ ) );
BUF_X1 \u0_ps2_kb/_0843_ ( .A(\u0_ps2_kb/_0151_ ), .Z(\u0_ps2_kb/_0055_ ) );
BUF_X1 \u0_ps2_kb/_0844_ ( .A(\u0_ps2_kb/fifo[4][2] ), .Z(\u0_ps2_kb/_0249_ ) );
BUF_X1 \u0_ps2_kb/_0845_ ( .A(\u0_ps2_kb/_0152_ ), .Z(\u0_ps2_kb/_0056_ ) );
BUF_X1 \u0_ps2_kb/_0846_ ( .A(\u0_ps2_kb/fifo[4][3] ), .Z(\u0_ps2_kb/_0250_ ) );
BUF_X1 \u0_ps2_kb/_0847_ ( .A(\u0_ps2_kb/_0153_ ), .Z(\u0_ps2_kb/_0057_ ) );
BUF_X1 \u0_ps2_kb/_0848_ ( .A(\u0_ps2_kb/fifo[4][4] ), .Z(\u0_ps2_kb/_0251_ ) );
BUF_X1 \u0_ps2_kb/_0849_ ( .A(\u0_ps2_kb/_0154_ ), .Z(\u0_ps2_kb/_0058_ ) );
BUF_X1 \u0_ps2_kb/_0850_ ( .A(\u0_ps2_kb/fifo[4][5] ), .Z(\u0_ps2_kb/_0252_ ) );
BUF_X1 \u0_ps2_kb/_0851_ ( .A(\u0_ps2_kb/_0155_ ), .Z(\u0_ps2_kb/_0059_ ) );
BUF_X1 \u0_ps2_kb/_0852_ ( .A(\u0_ps2_kb/fifo[4][6] ), .Z(\u0_ps2_kb/_0253_ ) );
BUF_X1 \u0_ps2_kb/_0853_ ( .A(\u0_ps2_kb/_0156_ ), .Z(\u0_ps2_kb/_0060_ ) );
BUF_X1 \u0_ps2_kb/_0854_ ( .A(\u0_ps2_kb/fifo[4][7] ), .Z(\u0_ps2_kb/_0254_ ) );
BUF_X1 \u0_ps2_kb/_0855_ ( .A(\u0_ps2_kb/_0157_ ), .Z(\u0_ps2_kb/_0061_ ) );
BUF_X1 \u0_ps2_kb/_0856_ ( .A(\u0_ps2_kb/fifo[0][0] ), .Z(\u0_ps2_kb/_0215_ ) );
BUF_X1 \u0_ps2_kb/_0857_ ( .A(\u0_ps2_kb/fifo[1][0] ), .Z(\u0_ps2_kb/_0223_ ) );
BUF_X1 \u0_ps2_kb/_0858_ ( .A(\u0_ps2_kb/r_ptr [0] ), .Z(\u0_ps2_kb/_0442_ ) );
BUF_X1 \u0_ps2_kb/_0859_ ( .A(\u0_ps2_kb/fifo[2][0] ), .Z(\u0_ps2_kb/_0231_ ) );
BUF_X1 \u0_ps2_kb/_0860_ ( .A(\u0_ps2_kb/fifo[3][0] ), .Z(\u0_ps2_kb/_0239_ ) );
BUF_X1 \u0_ps2_kb/_0861_ ( .A(\u0_ps2_kb/r_ptr [1] ), .Z(\u0_ps2_kb/_0443_ ) );
BUF_X1 \u0_ps2_kb/_0862_ ( .A(\u0_ps2_kb/fifo[5][0] ), .Z(\u0_ps2_kb/_0255_ ) );
BUF_X1 \u0_ps2_kb/_0863_ ( .A(\u0_ps2_kb/r_ptr [2] ), .Z(\u0_ps2_kb/_0444_ ) );
BUF_X1 \u0_ps2_kb/_0864_ ( .A(\u0_ps2_kb/_0207_ ), .Z(\data [0] ) );
BUF_X1 \u0_ps2_kb/_0865_ ( .A(\u0_ps2_kb/fifo[0][1] ), .Z(\u0_ps2_kb/_0216_ ) );
BUF_X1 \u0_ps2_kb/_0866_ ( .A(\u0_ps2_kb/fifo[1][1] ), .Z(\u0_ps2_kb/_0224_ ) );
BUF_X1 \u0_ps2_kb/_0867_ ( .A(\u0_ps2_kb/fifo[2][1] ), .Z(\u0_ps2_kb/_0232_ ) );
BUF_X1 \u0_ps2_kb/_0868_ ( .A(\u0_ps2_kb/fifo[3][1] ), .Z(\u0_ps2_kb/_0240_ ) );
BUF_X1 \u0_ps2_kb/_0869_ ( .A(\u0_ps2_kb/fifo[5][1] ), .Z(\u0_ps2_kb/_0256_ ) );
BUF_X1 \u0_ps2_kb/_0870_ ( .A(\u0_ps2_kb/_0208_ ), .Z(\data [1] ) );
BUF_X1 \u0_ps2_kb/_0871_ ( .A(\u0_ps2_kb/fifo[0][2] ), .Z(\u0_ps2_kb/_0217_ ) );
BUF_X1 \u0_ps2_kb/_0872_ ( .A(\u0_ps2_kb/fifo[1][2] ), .Z(\u0_ps2_kb/_0225_ ) );
BUF_X1 \u0_ps2_kb/_0873_ ( .A(\u0_ps2_kb/fifo[2][2] ), .Z(\u0_ps2_kb/_0233_ ) );
BUF_X1 \u0_ps2_kb/_0874_ ( .A(\u0_ps2_kb/fifo[3][2] ), .Z(\u0_ps2_kb/_0241_ ) );
BUF_X1 \u0_ps2_kb/_0875_ ( .A(\u0_ps2_kb/fifo[5][2] ), .Z(\u0_ps2_kb/_0257_ ) );
BUF_X1 \u0_ps2_kb/_0876_ ( .A(\u0_ps2_kb/_0209_ ), .Z(\data [2] ) );
BUF_X1 \u0_ps2_kb/_0877_ ( .A(\u0_ps2_kb/fifo[0][3] ), .Z(\u0_ps2_kb/_0218_ ) );
BUF_X1 \u0_ps2_kb/_0878_ ( .A(\u0_ps2_kb/fifo[1][3] ), .Z(\u0_ps2_kb/_0226_ ) );
BUF_X1 \u0_ps2_kb/_0879_ ( .A(\u0_ps2_kb/fifo[2][3] ), .Z(\u0_ps2_kb/_0234_ ) );
BUF_X1 \u0_ps2_kb/_0880_ ( .A(\u0_ps2_kb/fifo[3][3] ), .Z(\u0_ps2_kb/_0242_ ) );
BUF_X1 \u0_ps2_kb/_0881_ ( .A(\u0_ps2_kb/fifo[5][3] ), .Z(\u0_ps2_kb/_0258_ ) );
BUF_X1 \u0_ps2_kb/_0882_ ( .A(\u0_ps2_kb/_0210_ ), .Z(\data [3] ) );
BUF_X1 \u0_ps2_kb/_0883_ ( .A(\u0_ps2_kb/fifo[0][4] ), .Z(\u0_ps2_kb/_0219_ ) );
BUF_X1 \u0_ps2_kb/_0884_ ( .A(\u0_ps2_kb/fifo[1][4] ), .Z(\u0_ps2_kb/_0227_ ) );
BUF_X1 \u0_ps2_kb/_0885_ ( .A(\u0_ps2_kb/fifo[2][4] ), .Z(\u0_ps2_kb/_0235_ ) );
BUF_X1 \u0_ps2_kb/_0886_ ( .A(\u0_ps2_kb/fifo[3][4] ), .Z(\u0_ps2_kb/_0243_ ) );
BUF_X1 \u0_ps2_kb/_0887_ ( .A(\u0_ps2_kb/fifo[5][4] ), .Z(\u0_ps2_kb/_0259_ ) );
BUF_X1 \u0_ps2_kb/_0888_ ( .A(\u0_ps2_kb/_0211_ ), .Z(\data [4] ) );
BUF_X1 \u0_ps2_kb/_0889_ ( .A(\u0_ps2_kb/fifo[0][5] ), .Z(\u0_ps2_kb/_0220_ ) );
BUF_X1 \u0_ps2_kb/_0890_ ( .A(\u0_ps2_kb/fifo[1][5] ), .Z(\u0_ps2_kb/_0228_ ) );
BUF_X1 \u0_ps2_kb/_0891_ ( .A(\u0_ps2_kb/fifo[2][5] ), .Z(\u0_ps2_kb/_0236_ ) );
BUF_X1 \u0_ps2_kb/_0892_ ( .A(\u0_ps2_kb/fifo[3][5] ), .Z(\u0_ps2_kb/_0244_ ) );
BUF_X1 \u0_ps2_kb/_0893_ ( .A(\u0_ps2_kb/fifo[5][5] ), .Z(\u0_ps2_kb/_0260_ ) );
BUF_X1 \u0_ps2_kb/_0894_ ( .A(\u0_ps2_kb/_0212_ ), .Z(\data [5] ) );
BUF_X1 \u0_ps2_kb/_0895_ ( .A(\u0_ps2_kb/fifo[0][6] ), .Z(\u0_ps2_kb/_0221_ ) );
BUF_X1 \u0_ps2_kb/_0896_ ( .A(\u0_ps2_kb/fifo[1][6] ), .Z(\u0_ps2_kb/_0229_ ) );
BUF_X1 \u0_ps2_kb/_0897_ ( .A(\u0_ps2_kb/fifo[2][6] ), .Z(\u0_ps2_kb/_0237_ ) );
BUF_X1 \u0_ps2_kb/_0898_ ( .A(\u0_ps2_kb/fifo[3][6] ), .Z(\u0_ps2_kb/_0245_ ) );
BUF_X1 \u0_ps2_kb/_0899_ ( .A(\u0_ps2_kb/fifo[5][6] ), .Z(\u0_ps2_kb/_0261_ ) );
BUF_X1 \u0_ps2_kb/_0900_ ( .A(\u0_ps2_kb/_0213_ ), .Z(\data [6] ) );
BUF_X1 \u0_ps2_kb/_0901_ ( .A(\u0_ps2_kb/fifo[0][7] ), .Z(\u0_ps2_kb/_0222_ ) );
BUF_X1 \u0_ps2_kb/_0902_ ( .A(\u0_ps2_kb/fifo[1][7] ), .Z(\u0_ps2_kb/_0230_ ) );
BUF_X1 \u0_ps2_kb/_0903_ ( .A(\u0_ps2_kb/fifo[2][7] ), .Z(\u0_ps2_kb/_0238_ ) );
BUF_X1 \u0_ps2_kb/_0904_ ( .A(\u0_ps2_kb/fifo[3][7] ), .Z(\u0_ps2_kb/_0246_ ) );
BUF_X1 \u0_ps2_kb/_0905_ ( .A(\u0_ps2_kb/fifo[5][7] ), .Z(\u0_ps2_kb/_0262_ ) );
BUF_X1 \u0_ps2_kb/_0906_ ( .A(\u0_ps2_kb/_0214_ ), .Z(\data [7] ) );
BUF_X1 \u0_ps2_kb/_0907_ ( .A(\u0_ps2_kb/_0088_ ), .Z(\u0_ps2_kb/_0184_ ) );
BUF_X1 \u0_ps2_kb/_0908_ ( .A(\u0_ps2_kb/_0142_ ), .Z(\u0_ps2_kb/_0046_ ) );
BUF_X1 \u0_ps2_kb/_0909_ ( .A(\u0_ps2_kb/_0143_ ), .Z(\u0_ps2_kb/_0047_ ) );
BUF_X1 \u0_ps2_kb/_0910_ ( .A(\u0_ps2_kb/_0144_ ), .Z(\u0_ps2_kb/_0048_ ) );
BUF_X1 \u0_ps2_kb/_0911_ ( .A(\u0_ps2_kb/_0145_ ), .Z(\u0_ps2_kb/_0049_ ) );
BUF_X1 \u0_ps2_kb/_0912_ ( .A(\u0_ps2_kb/_0146_ ), .Z(\u0_ps2_kb/_0050_ ) );
BUF_X1 \u0_ps2_kb/_0913_ ( .A(\u0_ps2_kb/_0147_ ), .Z(\u0_ps2_kb/_0051_ ) );
BUF_X1 \u0_ps2_kb/_0914_ ( .A(\u0_ps2_kb/_0148_ ), .Z(\u0_ps2_kb/_0052_ ) );
BUF_X1 \u0_ps2_kb/_0915_ ( .A(\u0_ps2_kb/_0149_ ), .Z(\u0_ps2_kb/_0053_ ) );
BUF_X1 \u0_ps2_kb/_0916_ ( .A(\u0_ps2_kb/_0134_ ), .Z(\u0_ps2_kb/_0038_ ) );
BUF_X1 \u0_ps2_kb/_0917_ ( .A(\u0_ps2_kb/_0135_ ), .Z(\u0_ps2_kb/_0039_ ) );
BUF_X1 \u0_ps2_kb/_0918_ ( .A(\u0_ps2_kb/_0136_ ), .Z(\u0_ps2_kb/_0040_ ) );
BUF_X1 \u0_ps2_kb/_0919_ ( .A(\u0_ps2_kb/_0137_ ), .Z(\u0_ps2_kb/_0041_ ) );
BUF_X1 \u0_ps2_kb/_0920_ ( .A(\u0_ps2_kb/_0138_ ), .Z(\u0_ps2_kb/_0042_ ) );
BUF_X1 \u0_ps2_kb/_0921_ ( .A(\u0_ps2_kb/_0139_ ), .Z(\u0_ps2_kb/_0043_ ) );
BUF_X1 \u0_ps2_kb/_0922_ ( .A(\u0_ps2_kb/_0140_ ), .Z(\u0_ps2_kb/_0044_ ) );
BUF_X1 \u0_ps2_kb/_0923_ ( .A(\u0_ps2_kb/_0141_ ), .Z(\u0_ps2_kb/_0045_ ) );
BUF_X1 \u0_ps2_kb/_0924_ ( .A(\u0_ps2_kb/_0126_ ), .Z(\u0_ps2_kb/_0030_ ) );
BUF_X1 \u0_ps2_kb/_0925_ ( .A(\u0_ps2_kb/_0127_ ), .Z(\u0_ps2_kb/_0031_ ) );
BUF_X1 \u0_ps2_kb/_0926_ ( .A(\u0_ps2_kb/_0128_ ), .Z(\u0_ps2_kb/_0032_ ) );
BUF_X1 \u0_ps2_kb/_0927_ ( .A(\u0_ps2_kb/_0129_ ), .Z(\u0_ps2_kb/_0033_ ) );
BUF_X1 \u0_ps2_kb/_0928_ ( .A(\u0_ps2_kb/_0130_ ), .Z(\u0_ps2_kb/_0034_ ) );
BUF_X1 \u0_ps2_kb/_0929_ ( .A(\u0_ps2_kb/_0131_ ), .Z(\u0_ps2_kb/_0035_ ) );
BUF_X1 \u0_ps2_kb/_0930_ ( .A(\u0_ps2_kb/_0132_ ), .Z(\u0_ps2_kb/_0036_ ) );
BUF_X1 \u0_ps2_kb/_0931_ ( .A(\u0_ps2_kb/_0133_ ), .Z(\u0_ps2_kb/_0037_ ) );
BUF_X1 \u0_ps2_kb/_0932_ ( .A(\u0_ps2_kb/_0118_ ), .Z(\u0_ps2_kb/_0022_ ) );
BUF_X1 \u0_ps2_kb/_0933_ ( .A(\u0_ps2_kb/_0119_ ), .Z(\u0_ps2_kb/_0023_ ) );
BUF_X1 \u0_ps2_kb/_0934_ ( .A(\u0_ps2_kb/_0120_ ), .Z(\u0_ps2_kb/_0024_ ) );
BUF_X1 \u0_ps2_kb/_0935_ ( .A(\u0_ps2_kb/_0121_ ), .Z(\u0_ps2_kb/_0025_ ) );
BUF_X1 \u0_ps2_kb/_0936_ ( .A(\u0_ps2_kb/_0122_ ), .Z(\u0_ps2_kb/_0026_ ) );
BUF_X1 \u0_ps2_kb/_0937_ ( .A(\u0_ps2_kb/_0123_ ), .Z(\u0_ps2_kb/_0027_ ) );
BUF_X1 \u0_ps2_kb/_0938_ ( .A(\u0_ps2_kb/_0124_ ), .Z(\u0_ps2_kb/_0028_ ) );
BUF_X1 \u0_ps2_kb/_0939_ ( .A(\u0_ps2_kb/_0125_ ), .Z(\u0_ps2_kb/_0029_ ) );
BUF_X1 \u0_ps2_kb/_0940_ ( .A(\u0_ps2_kb/_0098_ ), .Z(\u0_ps2_kb/_0002_ ) );
BUF_X1 \u0_ps2_kb/_0941_ ( .A(\u0_ps2_kb/_0097_ ), .Z(\u0_ps2_kb/_0001_ ) );
BUF_X1 \u0_ps2_kb/_0942_ ( .A(\u0_ps2_kb/_0096_ ), .Z(\u0_ps2_kb/_0000_ ) );
BUF_X1 \u0_ps2_kb/_0943_ ( .A(\u0_ps2_kb/_0106_ ), .Z(\u0_ps2_kb/_0010_ ) );
BUF_X1 \u0_ps2_kb/_0944_ ( .A(\u0_ps2_kb/_0089_ ), .Z(\u0_ps2_kb/_0185_ ) );
BUF_X1 \u0_ps2_kb/_0945_ ( .A(\u0_ps2_kb/_0107_ ), .Z(\u0_ps2_kb/_0011_ ) );
BUF_X1 \u0_ps2_kb/_0946_ ( .A(\u0_ps2_kb/_0090_ ), .Z(\u0_ps2_kb/_0186_ ) );
BUF_X1 \u0_ps2_kb/_0947_ ( .A(\u0_ps2_kb/_0108_ ), .Z(\u0_ps2_kb/_0012_ ) );
BUF_X1 \u0_ps2_kb/_0948_ ( .A(\u0_ps2_kb/_0091_ ), .Z(\u0_ps2_kb/_0187_ ) );
BUF_X1 \u0_ps2_kb/_0949_ ( .A(\u0_ps2_kb/_0109_ ), .Z(\u0_ps2_kb/_0013_ ) );
BUF_X1 \u0_ps2_kb/_0950_ ( .A(nextdata_n ), .Z(\u0_ps2_kb/_0437_ ) );
BUF_X1 \u0_ps2_kb/_0951_ ( .A(\u0_ps2_kb/_0092_ ), .Z(\u0_ps2_kb/_0188_ ) );
BUF_X1 \u0_ps2_kb/_0952_ ( .A(ready ), .Z(\u0_ps2_kb/_0445_ ) );
BUF_X1 \u0_ps2_kb/_0953_ ( .A(\u0_ps2_kb/_0111_ ), .Z(\u0_ps2_kb/_0015_ ) );
BUF_X1 \u0_ps2_kb/_0954_ ( .A(\u0_ps2_kb/_0087_ ), .Z(\u0_ps2_kb/_0183_ ) );
BUF_X1 \u0_ps2_kb/_0955_ ( .A(\u0_ps2_kb/_0112_ ), .Z(\u0_ps2_kb/_0016_ ) );
BUF_X1 \u0_ps2_kb/_0956_ ( .A(\u0_ps2_kb/_0086_ ), .Z(\u0_ps2_kb/_0182_ ) );
BUF_X1 \u0_ps2_kb/_0957_ ( .A(\u0_ps2_kb/_0113_ ), .Z(\u0_ps2_kb/_0017_ ) );
BUF_X1 \u0_ps2_kb/_0958_ ( .A(\u0_ps2_kb/_0115_ ), .Z(\u0_ps2_kb/_0019_ ) );
BUF_X1 \u0_ps2_kb/_0959_ ( .A(\u0_ps2_kb/_0093_ ), .Z(\u0_ps2_kb/_0189_ ) );
BUF_X1 \u0_ps2_kb/_0960_ ( .A(\u0_ps2_kb/_0116_ ), .Z(\u0_ps2_kb/_0020_ ) );
BUF_X1 \u0_ps2_kb/_0961_ ( .A(\u0_ps2_kb/_0094_ ), .Z(\u0_ps2_kb/_0190_ ) );
BUF_X1 \u0_ps2_kb/_0962_ ( .A(\u0_ps2_kb/_0117_ ), .Z(\u0_ps2_kb/_0021_ ) );
BUF_X1 \u0_ps2_kb/_0963_ ( .A(\u0_ps2_kb/_0158_ ), .Z(\u0_ps2_kb/_0062_ ) );
BUF_X1 \u0_ps2_kb/_0964_ ( .A(\u0_ps2_kb/_0159_ ), .Z(\u0_ps2_kb/_0063_ ) );
BUF_X1 \u0_ps2_kb/_0965_ ( .A(\u0_ps2_kb/_0160_ ), .Z(\u0_ps2_kb/_0064_ ) );
BUF_X1 \u0_ps2_kb/_0966_ ( .A(\u0_ps2_kb/_0161_ ), .Z(\u0_ps2_kb/_0065_ ) );
BUF_X1 \u0_ps2_kb/_0967_ ( .A(\u0_ps2_kb/_0162_ ), .Z(\u0_ps2_kb/_0066_ ) );
BUF_X1 \u0_ps2_kb/_0968_ ( .A(\u0_ps2_kb/_0163_ ), .Z(\u0_ps2_kb/_0067_ ) );
BUF_X1 \u0_ps2_kb/_0969_ ( .A(\u0_ps2_kb/_0164_ ), .Z(\u0_ps2_kb/_0068_ ) );
BUF_X1 \u0_ps2_kb/_0970_ ( .A(\u0_ps2_kb/_0165_ ), .Z(\u0_ps2_kb/_0069_ ) );
BUF_X1 \u0_ps2_kb/_0971_ ( .A(\u0_ps2_kb/_0114_ ), .Z(\u0_ps2_kb/_0018_ ) );
BUF_X1 \u0_ps2_kb/_0972_ ( .A(overflow ), .Z(\u0_ps2_kb/_0438_ ) );
BUF_X1 \u0_ps2_kb/_0973_ ( .A(\u0_ps2_kb/_0095_ ), .Z(\u0_ps2_kb/_0191_ ) );
BUF_X1 \u0_ps2_kb/_0974_ ( .A(\u0_ps2_kb/_0110_ ), .Z(\u0_ps2_kb/_0014_ ) );
DFF_X1 \u0_ps2_kb/_0975_ ( .D(\u0_ps2_kb/_0070_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][0] ), .QN(\u0_ps2_kb/_0449_ ) );
DFF_X1 \u0_ps2_kb/_0976_ ( .D(\u0_ps2_kb/_0071_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][1] ), .QN(\u0_ps2_kb/_0450_ ) );
DFF_X1 \u0_ps2_kb/_0977_ ( .D(\u0_ps2_kb/_0072_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][2] ), .QN(\u0_ps2_kb/_0451_ ) );
DFF_X1 \u0_ps2_kb/_0978_ ( .D(\u0_ps2_kb/_0073_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][3] ), .QN(\u0_ps2_kb/_0452_ ) );
DFF_X1 \u0_ps2_kb/_0979_ ( .D(\u0_ps2_kb/_0074_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][4] ), .QN(\u0_ps2_kb/_0453_ ) );
DFF_X1 \u0_ps2_kb/_0980_ ( .D(\u0_ps2_kb/_0075_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][5] ), .QN(\u0_ps2_kb/_0454_ ) );
DFF_X1 \u0_ps2_kb/_0981_ ( .D(\u0_ps2_kb/_0076_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][6] ), .QN(\u0_ps2_kb/_0455_ ) );
DFF_X1 \u0_ps2_kb/_0982_ ( .D(\u0_ps2_kb/_0077_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][7] ), .QN(\u0_ps2_kb/_0456_ ) );
DFF_X1 \u0_ps2_kb/_0983_ ( .D(\u0_ps2_kb/_0062_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][0] ), .QN(\u0_ps2_kb/_0457_ ) );
DFF_X1 \u0_ps2_kb/_0984_ ( .D(\u0_ps2_kb/_0063_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][1] ), .QN(\u0_ps2_kb/_0458_ ) );
DFF_X1 \u0_ps2_kb/_0985_ ( .D(\u0_ps2_kb/_0064_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][2] ), .QN(\u0_ps2_kb/_0459_ ) );
DFF_X1 \u0_ps2_kb/_0986_ ( .D(\u0_ps2_kb/_0065_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][3] ), .QN(\u0_ps2_kb/_0460_ ) );
DFF_X1 \u0_ps2_kb/_0987_ ( .D(\u0_ps2_kb/_0066_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][4] ), .QN(\u0_ps2_kb/_0461_ ) );
DFF_X1 \u0_ps2_kb/_0988_ ( .D(\u0_ps2_kb/_0067_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][5] ), .QN(\u0_ps2_kb/_0462_ ) );
DFF_X1 \u0_ps2_kb/_0989_ ( .D(\u0_ps2_kb/_0068_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][6] ), .QN(\u0_ps2_kb/_0463_ ) );
DFF_X1 \u0_ps2_kb/_0990_ ( .D(\u0_ps2_kb/_0069_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][7] ), .QN(\u0_ps2_kb/_0464_ ) );
DFF_X1 \u0_ps2_kb/_0991_ ( .D(\u0_ps2_kb/_0015_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr [0] ), .QN(\u0_ps2_kb/_0092_ ) );
DFF_X1 \u0_ps2_kb/_0992_ ( .D(\u0_ps2_kb/_0016_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr [1] ), .QN(\u0_ps2_kb/_0087_ ) );
DFF_X1 \u0_ps2_kb/_0993_ ( .D(\u0_ps2_kb/_0017_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr [2] ), .QN(\u0_ps2_kb/_0086_ ) );
DFF_X1 \u0_ps2_kb/_0994_ ( .D(\u0_ps2_kb/_0078_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][0] ), .QN(\u0_ps2_kb/_0465_ ) );
DFF_X1 \u0_ps2_kb/_0995_ ( .D(\u0_ps2_kb/_0079_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][1] ), .QN(\u0_ps2_kb/_0466_ ) );
DFF_X1 \u0_ps2_kb/_0996_ ( .D(\u0_ps2_kb/_0080_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][2] ), .QN(\u0_ps2_kb/_0467_ ) );
DFF_X1 \u0_ps2_kb/_0997_ ( .D(\u0_ps2_kb/_0081_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][3] ), .QN(\u0_ps2_kb/_0468_ ) );
DFF_X1 \u0_ps2_kb/_0998_ ( .D(\u0_ps2_kb/_0082_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][4] ), .QN(\u0_ps2_kb/_0469_ ) );
DFF_X1 \u0_ps2_kb/_0999_ ( .D(\u0_ps2_kb/_0083_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][5] ), .QN(\u0_ps2_kb/_0470_ ) );
DFF_X1 \u0_ps2_kb/_1000_ ( .D(\u0_ps2_kb/_0084_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][6] ), .QN(\u0_ps2_kb/_0471_ ) );
DFF_X1 \u0_ps2_kb/_1001_ ( .D(\u0_ps2_kb/_0085_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][7] ), .QN(\u0_ps2_kb/_0472_ ) );
DFF_X1 \u0_ps2_kb/_1002_ ( .D(\u0_ps2_kb/_0022_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][0] ), .QN(\u0_ps2_kb/_0473_ ) );
DFF_X1 \u0_ps2_kb/_1003_ ( .D(\u0_ps2_kb/_0023_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][1] ), .QN(\u0_ps2_kb/_0474_ ) );
DFF_X1 \u0_ps2_kb/_1004_ ( .D(\u0_ps2_kb/_0024_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][2] ), .QN(\u0_ps2_kb/_0475_ ) );
DFF_X1 \u0_ps2_kb/_1005_ ( .D(\u0_ps2_kb/_0025_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][3] ), .QN(\u0_ps2_kb/_0476_ ) );
DFF_X1 \u0_ps2_kb/_1006_ ( .D(\u0_ps2_kb/_0026_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][4] ), .QN(\u0_ps2_kb/_0477_ ) );
DFF_X1 \u0_ps2_kb/_1007_ ( .D(\u0_ps2_kb/_0027_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][5] ), .QN(\u0_ps2_kb/_0478_ ) );
DFF_X1 \u0_ps2_kb/_1008_ ( .D(\u0_ps2_kb/_0028_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][6] ), .QN(\u0_ps2_kb/_0479_ ) );
DFF_X1 \u0_ps2_kb/_1009_ ( .D(\u0_ps2_kb/_0029_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][7] ), .QN(\u0_ps2_kb/_0480_ ) );
DFF_X1 \u0_ps2_kb/_1010_ ( .D(\u0_ps2_kb/_0046_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][0] ), .QN(\u0_ps2_kb/_0481_ ) );
DFF_X1 \u0_ps2_kb/_1011_ ( .D(\u0_ps2_kb/_0047_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][1] ), .QN(\u0_ps2_kb/_0482_ ) );
DFF_X1 \u0_ps2_kb/_1012_ ( .D(\u0_ps2_kb/_0048_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][2] ), .QN(\u0_ps2_kb/_0483_ ) );
DFF_X1 \u0_ps2_kb/_1013_ ( .D(\u0_ps2_kb/_0049_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][3] ), .QN(\u0_ps2_kb/_0484_ ) );
DFF_X1 \u0_ps2_kb/_1014_ ( .D(\u0_ps2_kb/_0050_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][4] ), .QN(\u0_ps2_kb/_0485_ ) );
DFF_X1 \u0_ps2_kb/_1015_ ( .D(\u0_ps2_kb/_0051_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][5] ), .QN(\u0_ps2_kb/_0486_ ) );
DFF_X1 \u0_ps2_kb/_1016_ ( .D(\u0_ps2_kb/_0052_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][6] ), .QN(\u0_ps2_kb/_0487_ ) );
DFF_X1 \u0_ps2_kb/_1017_ ( .D(\u0_ps2_kb/_0053_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][7] ), .QN(\u0_ps2_kb/_0488_ ) );
DFF_X1 \u0_ps2_kb/_1018_ ( .D(\u0_ps2_kb/_0054_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][0] ), .QN(\u0_ps2_kb/_0489_ ) );
DFF_X1 \u0_ps2_kb/_1019_ ( .D(\u0_ps2_kb/_0055_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][1] ), .QN(\u0_ps2_kb/_0490_ ) );
DFF_X1 \u0_ps2_kb/_1020_ ( .D(\u0_ps2_kb/_0056_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][2] ), .QN(\u0_ps2_kb/_0491_ ) );
DFF_X1 \u0_ps2_kb/_1021_ ( .D(\u0_ps2_kb/_0057_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][3] ), .QN(\u0_ps2_kb/_0492_ ) );
DFF_X1 \u0_ps2_kb/_1022_ ( .D(\u0_ps2_kb/_0058_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][4] ), .QN(\u0_ps2_kb/_0493_ ) );
DFF_X1 \u0_ps2_kb/_1023_ ( .D(\u0_ps2_kb/_0059_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][5] ), .QN(\u0_ps2_kb/_0494_ ) );
DFF_X1 \u0_ps2_kb/_1024_ ( .D(\u0_ps2_kb/_0060_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][6] ), .QN(\u0_ps2_kb/_0495_ ) );
DFF_X1 \u0_ps2_kb/_1025_ ( .D(\u0_ps2_kb/_0061_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][7] ), .QN(\u0_ps2_kb/_0496_ ) );
DFF_X1 \u0_ps2_kb/_1026_ ( .D(\u0_ps2_kb/_0038_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][0] ), .QN(\u0_ps2_kb/_0497_ ) );
DFF_X1 \u0_ps2_kb/_1027_ ( .D(\u0_ps2_kb/_0039_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][1] ), .QN(\u0_ps2_kb/_0498_ ) );
DFF_X1 \u0_ps2_kb/_1028_ ( .D(\u0_ps2_kb/_0040_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][2] ), .QN(\u0_ps2_kb/_0499_ ) );
DFF_X1 \u0_ps2_kb/_1029_ ( .D(\u0_ps2_kb/_0041_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][3] ), .QN(\u0_ps2_kb/_0500_ ) );
DFF_X1 \u0_ps2_kb/_1030_ ( .D(\u0_ps2_kb/_0042_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][4] ), .QN(\u0_ps2_kb/_0501_ ) );
DFF_X1 \u0_ps2_kb/_1031_ ( .D(\u0_ps2_kb/_0043_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][5] ), .QN(\u0_ps2_kb/_0502_ ) );
DFF_X1 \u0_ps2_kb/_1032_ ( .D(\u0_ps2_kb/_0044_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][6] ), .QN(\u0_ps2_kb/_0503_ ) );
DFF_X1 \u0_ps2_kb/_1033_ ( .D(\u0_ps2_kb/_0045_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][7] ), .QN(\u0_ps2_kb/_0504_ ) );
DFF_X1 \u0_ps2_kb/_1034_ ( .D(\u0_ps2_kb/_0030_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][0] ), .QN(\u0_ps2_kb/_0505_ ) );
DFF_X1 \u0_ps2_kb/_1035_ ( .D(\u0_ps2_kb/_0031_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][1] ), .QN(\u0_ps2_kb/_0506_ ) );
DFF_X1 \u0_ps2_kb/_1036_ ( .D(\u0_ps2_kb/_0032_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][2] ), .QN(\u0_ps2_kb/_0507_ ) );
DFF_X1 \u0_ps2_kb/_1037_ ( .D(\u0_ps2_kb/_0033_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][3] ), .QN(\u0_ps2_kb/_0508_ ) );
DFF_X1 \u0_ps2_kb/_1038_ ( .D(\u0_ps2_kb/_0034_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][4] ), .QN(\u0_ps2_kb/_0509_ ) );
DFF_X1 \u0_ps2_kb/_1039_ ( .D(\u0_ps2_kb/_0035_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][5] ), .QN(\u0_ps2_kb/_0510_ ) );
DFF_X1 \u0_ps2_kb/_1040_ ( .D(\u0_ps2_kb/_0036_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][6] ), .QN(\u0_ps2_kb/_0511_ ) );
DFF_X1 \u0_ps2_kb/_1041_ ( .D(\u0_ps2_kb/_0037_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][7] ), .QN(\u0_ps2_kb/_0512_ ) );
DFF_X1 \u0_ps2_kb/_1042_ ( .D(\u0_ps2_kb/_0014_ ), .CK(clk ), .Q(overflow ), .QN(\u0_ps2_kb/_0095_ ) );
DFF_X1 \u0_ps2_kb/_1043_ ( .D(\u0_ps2_kb/_0018_ ), .CK(clk ), .Q(ready ), .QN(\u0_ps2_kb/_0513_ ) );
DFF_X1 \u0_ps2_kb/_1044_ ( .D(\u0_ps2_kb/_0000_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [0] ), .QN(\u0_ps2_kb/_0514_ ) );
DFF_X1 \u0_ps2_kb/_1045_ ( .D(\u0_ps2_kb/_0001_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [1] ), .QN(\u0_ps2_kb/_0515_ ) );
DFF_X1 \u0_ps2_kb/_1046_ ( .D(\u0_ps2_kb/_0002_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [2] ), .QN(\u0_ps2_kb/_0516_ ) );
DFF_X1 \u0_ps2_kb/_1047_ ( .D(\u0_ps2_kb/_0003_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [3] ), .QN(\u0_ps2_kb/_0517_ ) );
DFF_X1 \u0_ps2_kb/_1048_ ( .D(\u0_ps2_kb/_0004_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [4] ), .QN(\u0_ps2_kb/_0518_ ) );
DFF_X1 \u0_ps2_kb/_1049_ ( .D(\u0_ps2_kb/_0005_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [5] ), .QN(\u0_ps2_kb/_0519_ ) );
DFF_X1 \u0_ps2_kb/_1050_ ( .D(\u0_ps2_kb/_0006_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [6] ), .QN(\u0_ps2_kb/_0520_ ) );
DFF_X1 \u0_ps2_kb/_1051_ ( .D(\u0_ps2_kb/_0007_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [7] ), .QN(\u0_ps2_kb/_0521_ ) );
DFF_X1 \u0_ps2_kb/_1052_ ( .D(\u0_ps2_kb/_0008_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [8] ), .QN(\u0_ps2_kb/_0522_ ) );
DFF_X1 \u0_ps2_kb/_1053_ ( .D(\u0_ps2_kb/_0009_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer [9] ), .QN(\u0_ps2_kb/_0523_ ) );
DFF_X1 \u0_ps2_kb/_1054_ ( .D(\u0_ps2_kb/_0019_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr [0] ), .QN(\u0_ps2_kb/_0088_ ) );
DFF_X1 \u0_ps2_kb/_1055_ ( .D(\u0_ps2_kb/_0020_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr [1] ), .QN(\u0_ps2_kb/_0093_ ) );
DFF_X1 \u0_ps2_kb/_1056_ ( .D(\u0_ps2_kb/_0021_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr [2] ), .QN(\u0_ps2_kb/_0094_ ) );
DFF_X1 \u0_ps2_kb/_1057_ ( .D(\u0_ps2_kb/_0010_ ), .CK(clk ), .Q(\u0_ps2_kb/count [0] ), .QN(\u0_ps2_kb/_0524_ ) );
DFF_X1 \u0_ps2_kb/_1058_ ( .D(\u0_ps2_kb/_0011_ ), .CK(clk ), .Q(\u0_ps2_kb/count [1] ), .QN(\u0_ps2_kb/_0089_ ) );
DFF_X1 \u0_ps2_kb/_1059_ ( .D(\u0_ps2_kb/_0012_ ), .CK(clk ), .Q(\u0_ps2_kb/count [2] ), .QN(\u0_ps2_kb/_0090_ ) );
DFF_X1 \u0_ps2_kb/_1060_ ( .D(\u0_ps2_kb/_0013_ ), .CK(clk ), .Q(\u0_ps2_kb/count [3] ), .QN(\u0_ps2_kb/_0091_ ) );
DFF_X1 \u0_ps2_kb/_1061_ ( .D(ps2_clk ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync [0] ), .QN(\u0_ps2_kb/_0525_ ) );
DFF_X1 \u0_ps2_kb/_1062_ ( .D(\u0_ps2_kb/ps2_clk_sync [0] ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync [1] ), .QN(\u0_ps2_kb/_0526_ ) );
DFF_X1 \u0_ps2_kb/_1063_ ( .D(\u0_ps2_kb/ps2_clk_sync [1] ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync [2] ), .QN(\u0_ps2_kb/_0527_ ) );
NOR4_X2 \u1_ps2_dsh/_052_ ( .A1(\u1_ps2_dsh/_027_ ), .A2(\u1_ps2_dsh/_026_ ), .A3(\u1_ps2_dsh/_029_ ), .A4(\u1_ps2_dsh/_028_ ), .ZN(\u1_ps2_dsh/_034_ ) );
AND4_X1 \u1_ps2_dsh/_053_ ( .A1(\u1_ps2_dsh/_031_ ), .A2(\u1_ps2_dsh/_030_ ), .A3(\u1_ps2_dsh/_033_ ), .A4(\u1_ps2_dsh/_032_ ), .ZN(\u1_ps2_dsh/_035_ ) );
AND2_X1 \u1_ps2_dsh/_054_ ( .A1(\u1_ps2_dsh/_034_ ), .A2(\u1_ps2_dsh/_035_ ), .ZN(\u1_ps2_dsh/_017_ ) );
NAND2_X1 \u1_ps2_dsh/_055_ ( .A1(\u1_ps2_dsh/_031_ ), .A2(\u1_ps2_dsh/_032_ ), .ZN(\u1_ps2_dsh/_036_ ) );
NOR3_X2 \u1_ps2_dsh/_056_ ( .A1(\u1_ps2_dsh/_036_ ), .A2(\u1_ps2_dsh/_026_ ), .A3(\u1_ps2_dsh/_029_ ), .ZN(\u1_ps2_dsh/_037_ ) );
NAND2_X1 \u1_ps2_dsh/_057_ ( .A1(\u1_ps2_dsh/_030_ ), .A2(\u1_ps2_dsh/_033_ ), .ZN(\u1_ps2_dsh/_038_ ) );
NOR3_X2 \u1_ps2_dsh/_058_ ( .A1(\u1_ps2_dsh/_038_ ), .A2(\u1_ps2_dsh/_027_ ), .A3(\u1_ps2_dsh/_028_ ), .ZN(\u1_ps2_dsh/_039_ ) );
NAND2_X2 \u1_ps2_dsh/_059_ ( .A1(\u1_ps2_dsh/_037_ ), .A2(\u1_ps2_dsh/_039_ ), .ZN(\u1_ps2_dsh/_040_ ) );
AND2_X1 \u1_ps2_dsh/_060_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_018_ ), .ZN(\u1_ps2_dsh/_009_ ) );
AND2_X1 \u1_ps2_dsh/_061_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_019_ ), .ZN(\u1_ps2_dsh/_010_ ) );
AND2_X1 \u1_ps2_dsh/_062_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_020_ ), .ZN(\u1_ps2_dsh/_011_ ) );
AND2_X1 \u1_ps2_dsh/_063_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_021_ ), .ZN(\u1_ps2_dsh/_012_ ) );
AND2_X1 \u1_ps2_dsh/_064_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_022_ ), .ZN(\u1_ps2_dsh/_013_ ) );
AND2_X1 \u1_ps2_dsh/_065_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_023_ ), .ZN(\u1_ps2_dsh/_014_ ) );
AND2_X1 \u1_ps2_dsh/_066_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_024_ ), .ZN(\u1_ps2_dsh/_015_ ) );
AND2_X1 \u1_ps2_dsh/_067_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_025_ ), .ZN(\u1_ps2_dsh/_016_ ) );
LOGIC1_X1 \u1_ps2_dsh/_068_ ( .Z(\u1_ps2_dsh/_050_ ) );
LOGIC0_X1 \u1_ps2_dsh/_069_ ( .Z(\u1_ps2_dsh/_051_ ) );
BUF_X1 \u1_ps2_dsh/_070_ ( .A(\data_d1 [1] ), .Z(\u1_ps2_dsh/_027_ ) );
BUF_X1 \u1_ps2_dsh/_071_ ( .A(\data_d1 [0] ), .Z(\u1_ps2_dsh/_026_ ) );
BUF_X1 \u1_ps2_dsh/_072_ ( .A(\data_d1 [3] ), .Z(\u1_ps2_dsh/_029_ ) );
BUF_X1 \u1_ps2_dsh/_073_ ( .A(\data_d1 [2] ), .Z(\u1_ps2_dsh/_028_ ) );
BUF_X1 \u1_ps2_dsh/_074_ ( .A(\data_d1 [5] ), .Z(\u1_ps2_dsh/_031_ ) );
BUF_X1 \u1_ps2_dsh/_075_ ( .A(\data_d1 [4] ), .Z(\u1_ps2_dsh/_030_ ) );
BUF_X1 \u1_ps2_dsh/_076_ ( .A(\data_d1 [7] ), .Z(\u1_ps2_dsh/_033_ ) );
BUF_X1 \u1_ps2_dsh/_077_ ( .A(\data_d1 [6] ), .Z(\u1_ps2_dsh/_032_ ) );
BUF_X1 \u1_ps2_dsh/_078_ ( .A(\u1_ps2_dsh/_017_ ), .Z(\u1_ps2_dsh/_008_ ) );
BUF_X1 \u1_ps2_dsh/_079_ ( .A(\u1_ps2_dsh/ascii_result [0] ), .Z(\u1_ps2_dsh/_018_ ) );
BUF_X1 \u1_ps2_dsh/_080_ ( .A(\u1_ps2_dsh/_009_ ), .Z(\u1_ps2_dsh/_000_ ) );
BUF_X1 \u1_ps2_dsh/_081_ ( .A(\u1_ps2_dsh/ascii_result [1] ), .Z(\u1_ps2_dsh/_019_ ) );
BUF_X1 \u1_ps2_dsh/_082_ ( .A(\u1_ps2_dsh/_010_ ), .Z(\u1_ps2_dsh/_001_ ) );
BUF_X1 \u1_ps2_dsh/_083_ ( .A(\u1_ps2_dsh/ascii_result [2] ), .Z(\u1_ps2_dsh/_020_ ) );
BUF_X1 \u1_ps2_dsh/_084_ ( .A(\u1_ps2_dsh/_011_ ), .Z(\u1_ps2_dsh/_002_ ) );
BUF_X1 \u1_ps2_dsh/_085_ ( .A(\u1_ps2_dsh/ascii_result [3] ), .Z(\u1_ps2_dsh/_021_ ) );
BUF_X1 \u1_ps2_dsh/_086_ ( .A(\u1_ps2_dsh/_012_ ), .Z(\u1_ps2_dsh/_003_ ) );
BUF_X1 \u1_ps2_dsh/_087_ ( .A(\u1_ps2_dsh/ascii_result [4] ), .Z(\u1_ps2_dsh/_022_ ) );
BUF_X1 \u1_ps2_dsh/_088_ ( .A(\u1_ps2_dsh/_013_ ), .Z(\u1_ps2_dsh/_004_ ) );
BUF_X1 \u1_ps2_dsh/_089_ ( .A(\u1_ps2_dsh/ascii_result [5] ), .Z(\u1_ps2_dsh/_023_ ) );
BUF_X1 \u1_ps2_dsh/_090_ ( .A(\u1_ps2_dsh/_014_ ), .Z(\u1_ps2_dsh/_005_ ) );
BUF_X1 \u1_ps2_dsh/_091_ ( .A(\u1_ps2_dsh/ascii_result [6] ), .Z(\u1_ps2_dsh/_024_ ) );
BUF_X1 \u1_ps2_dsh/_092_ ( .A(\u1_ps2_dsh/_015_ ), .Z(\u1_ps2_dsh/_006_ ) );
BUF_X1 \u1_ps2_dsh/_093_ ( .A(\u1_ps2_dsh/ascii_result [7] ), .Z(\u1_ps2_dsh/_025_ ) );
BUF_X1 \u1_ps2_dsh/_094_ ( .A(\u1_ps2_dsh/_016_ ), .Z(\u1_ps2_dsh/_007_ ) );
DFFR_X1 \u1_ps2_dsh/_095_ ( .D(\u1_ps2_dsh/_008_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(key_release ), .QN(\u1_ps2_dsh/_041_ ) );
DFFR_X1 \u1_ps2_dsh/_096_ ( .D(\u1_ps2_dsh/_000_ ), .RN(fanout_net_28 ), .CK(clk ), .Q(\ascii [0] ), .QN(\u1_ps2_dsh/_042_ ) );
DFFR_X1 \u1_ps2_dsh/_097_ ( .D(\u1_ps2_dsh/_001_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [1] ), .QN(\u1_ps2_dsh/_043_ ) );
DFFR_X1 \u1_ps2_dsh/_098_ ( .D(\u1_ps2_dsh/_002_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [2] ), .QN(\u1_ps2_dsh/_044_ ) );
DFFR_X1 \u1_ps2_dsh/_099_ ( .D(\u1_ps2_dsh/_003_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [3] ), .QN(\u1_ps2_dsh/_045_ ) );
DFFR_X1 \u1_ps2_dsh/_100_ ( .D(\u1_ps2_dsh/_004_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [4] ), .QN(\u1_ps2_dsh/_046_ ) );
DFFR_X1 \u1_ps2_dsh/_101_ ( .D(\u1_ps2_dsh/_005_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [5] ), .QN(\u1_ps2_dsh/_047_ ) );
DFFR_X1 \u1_ps2_dsh/_102_ ( .D(\u1_ps2_dsh/_006_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [6] ), .QN(\u1_ps2_dsh/_048_ ) );
DFFR_X1 \u1_ps2_dsh/_103_ ( .D(\u1_ps2_dsh/_007_ ), .RN(clrn ), .CK(clk ), .Q(\ascii [7] ), .QN(\u1_ps2_dsh/_049_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1344_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0450_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0937_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1345_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0449_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0938_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1346_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0454_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0939_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1347_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0453_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0940_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1348_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0937_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0938_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0939_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0940_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0941_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1349_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0446_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0942_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1350_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0451_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0943_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1351_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0447_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0944_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1352_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0452_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0945_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1353_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0942_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0943_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0944_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0945_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0946_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1354_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0947_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1355_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0551_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0948_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1356_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0550_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0949_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1357_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0546_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0950_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1358_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0545_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0951_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1359_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0948_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0949_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0950_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0951_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0952_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1360_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0548_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0953_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1361_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0537_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0954_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1362_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0549_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0955_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1363_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0544_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0956_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1364_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0953_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0954_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0955_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0956_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0957_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1365_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0958_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1366_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0486_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0959_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1367_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0485_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0960_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1368_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0490_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0961_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1369_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0489_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0962_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1370_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0959_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0960_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0961_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0962_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0963_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1371_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0483_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0964_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1372_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0487_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0965_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1373_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0484_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0966_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1374_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0488_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0967_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1375_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0964_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0965_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0966_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0967_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0968_ ) );
AND2_X2 \u1_ps2_dsh/key_ascii/i0/_1376_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0969_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1377_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0236_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0970_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1378_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0235_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0971_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1379_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0242_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0972_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1380_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0241_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0973_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1381_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0970_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0971_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0972_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0973_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0974_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1382_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0233_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0975_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1383_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0239_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0976_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1384_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0234_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0977_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1385_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0240_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0978_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1386_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0975_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0976_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0977_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0978_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0979_ ) );
AND2_X4 \u1_ps2_dsh/key_ascii/i0/_1387_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0980_ ) );
OR4_X4 \u1_ps2_dsh/key_ascii/i0/_1388_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0947_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0958_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0969_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0980_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0981_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1389_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0414_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0982_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1390_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0413_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0983_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1391_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0419_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0984_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1392_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0418_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0985_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1393_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0982_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0983_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0984_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0985_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0986_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1394_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0411_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0987_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1395_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0416_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0988_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1396_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0412_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0989_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1397_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0417_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0990_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1398_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0987_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0988_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0989_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0990_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0991_ ) );
AND2_X4 \u1_ps2_dsh/key_ascii/i0/_1399_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0986_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0991_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0992_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1400_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0131_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0993_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1401_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0130_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0994_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1402_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0135_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0995_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1403_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0134_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0996_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1404_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0993_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0994_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0995_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0996_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0997_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1405_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0128_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0998_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1406_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0132_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0999_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1407_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0129_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1000_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1408_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0133_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1001_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1409_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0998_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0999_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1000_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1001_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1002_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1410_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1003_ ) );
OR2_X1 \u1_ps2_dsh/key_ascii/i0/_1411_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0992_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1003_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1004_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1412_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0379_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1005_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1413_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0378_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1006_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1414_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0376_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1007_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1415_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0377_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1008_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1416_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1005_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1006_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1007_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1008_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1009_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1417_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0384_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1010_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1418_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0383_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1011_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1419_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0380_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1012_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1420_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0381_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1013_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1421_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1010_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1011_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1012_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1013_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1014_ ) );
NOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1422_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1009_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1014_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1015_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1423_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0166_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1016_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1424_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0165_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1017_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1425_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0170_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1018_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1426_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0169_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1019_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1427_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1016_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1017_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1018_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1019_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1020_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1428_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0163_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1021_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1429_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0167_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1022_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1430_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0164_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1023_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1431_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0168_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1024_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1432_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1021_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1022_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1023_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1024_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1025_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1433_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1026_ ) );
NOR4_X4 \u1_ps2_dsh/key_ascii/i0/_1434_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0981_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1004_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1026_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1027_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1435_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0223_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1028_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1436_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0222_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1029_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1437_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0219_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1030_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1438_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0218_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1031_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1439_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1028_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1029_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1030_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1031_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1032_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1440_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0220_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1033_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1441_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0216_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1034_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1442_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0221_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1035_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1443_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0217_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1036_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1444_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1033_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1034_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1035_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1036_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1037_ ) );
AND2_X2 \u1_ps2_dsh/key_ascii/i0/_1445_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1038_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1446_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0188_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1039_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1447_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0187_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1040_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1448_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0184_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1041_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1449_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0183_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1042_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1450_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1039_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1040_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1041_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1042_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1043_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1451_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0185_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1044_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1452_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0180_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1045_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1453_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0186_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1046_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1454_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0181_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1047_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1455_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1044_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1045_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1046_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1047_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1048_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1456_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1038_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1049_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1457_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0473_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1050_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1458_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0472_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1051_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1459_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0468_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1052_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1460_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0467_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1053_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1461_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1050_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1051_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1052_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1053_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1054_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1462_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0469_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1055_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1463_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0465_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1056_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1464_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0470_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1057_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1465_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0466_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1058_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1466_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1055_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1056_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1057_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1058_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1059_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1467_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0259_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1060_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1468_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0258_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1061_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1469_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0255_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1062_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1470_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0254_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1063_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1471_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1060_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1061_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1062_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1063_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1064_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1472_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0256_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1065_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1473_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0252_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1066_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1474_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0257_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1067_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1475_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0253_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1068_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1476_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1065_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1066_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1067_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1068_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1069_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1477_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1070_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1478_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0508_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1071_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1479_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0507_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1072_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1480_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0503_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1073_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1481_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0502_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1074_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1482_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1071_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1072_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1073_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1074_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1075_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1483_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0505_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1076_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1484_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0500_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1077_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1485_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0506_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1078_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1486_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0501_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1079_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1487_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1076_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1077_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1078_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1079_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1080_ ) );
NOR2_X4 \u1_ps2_dsh/key_ascii/i0/_1488_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1075_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1080_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1081_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1489_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0201_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1082_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1490_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0200_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1083_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1491_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0206_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1084_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1492_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0205_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1085_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1493_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1082_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1083_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1084_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1085_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1086_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1494_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0198_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1087_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1495_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1088_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1496_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0199_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1089_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1497_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0203_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1090_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1498_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1087_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1088_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1089_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1090_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1091_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1499_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1092_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1500_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0153_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1093_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1501_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0152_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1094_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1502_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0148_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1095_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1503_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0147_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1096_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1504_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1093_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1094_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1095_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1096_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1097_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1505_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0150_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1098_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1506_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0145_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1099_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1507_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0151_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1100_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1508_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0146_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1101_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1509_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1098_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1099_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1100_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1101_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1102_ ) );
NOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1510_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1097_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1102_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1103_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1511_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0543_ ), .B(fanout_net_27 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1104_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1512_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0542_ ), .B(fanout_net_26 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1105_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1513_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0539_ ), .B(fanout_net_23 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1106_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1514_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0538_ ), .B(fanout_net_22 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1107_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1515_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1104_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1105_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1106_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1107_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1108_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1516_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0540_ ), .B(fanout_net_24 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1109_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1517_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0535_ ), .B(fanout_net_20 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1110_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1518_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0541_ ), .B(fanout_net_25 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1111_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1519_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0536_ ), .B(fanout_net_21 ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1112_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1520_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1109_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1110_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1111_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1112_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1113_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1521_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1114_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1522_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1049_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1070_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1092_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1114_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1115_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1523_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0081_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1116_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1524_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0080_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1117_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1525_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0077_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1118_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1526_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0076_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1119_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1527_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1116_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1117_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1118_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1119_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1120_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1528_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0078_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1121_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1529_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0074_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1122_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1530_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0079_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1123_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1531_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0075_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1124_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1532_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1121_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1122_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1123_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1124_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1125_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1533_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0564_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1126_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1534_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0563_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1127_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1535_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0568_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1128_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1536_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0567_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1129_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1537_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1126_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1127_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1128_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1129_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1130_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1538_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0561_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1131_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1539_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0565_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1132_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1540_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0562_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1133_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1541_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0566_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1134_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1542_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1131_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1132_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1133_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1134_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1135_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1543_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1136_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1544_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0046_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1137_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1545_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0045_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1138_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1546_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0042_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1139_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1547_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0041_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1140_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1548_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1137_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1138_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1139_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1140_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1141_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1549_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0043_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1142_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1550_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0039_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1143_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1551_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0044_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1144_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1552_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0040_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1145_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1553_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1142_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1143_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1144_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1145_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1146_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1554_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0393_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1147_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1555_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0382_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1148_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1556_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0437_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1149_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1557_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0426_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1150_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1558_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1147_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1148_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1149_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1150_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1151_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1559_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0360_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1152_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1560_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0404_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1153_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1561_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0371_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1154_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1562_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0415_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1155_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1563_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1152_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1153_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1154_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1155_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1156_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1564_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1157_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1565_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1136_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1157_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1158_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1566_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0024_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1159_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1567_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0023_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1160_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1568_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0029_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1161_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1569_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0028_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1162_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1570_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1159_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1160_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1161_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1162_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1163_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1571_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0021_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1164_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1572_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0025_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1165_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1573_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0022_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1166_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1574_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0026_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1167_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1575_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1164_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1165_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1166_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1167_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1168_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1576_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1169_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1577_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0095_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1170_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1578_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0094_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1171_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1579_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0099_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1172_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1580_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0098_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1173_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1581_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1170_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1171_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1172_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1173_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1174_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1582_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0091_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1175_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1583_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0096_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1176_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1584_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0092_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1177_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1585_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0097_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1178_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1586_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1175_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1176_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1177_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1178_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1179_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1587_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1180_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1588_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0059_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1181_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1589_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0058_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1182_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1590_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0056_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1183_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1591_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0057_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1184_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1592_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1181_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1182_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1183_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1184_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1185_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1593_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0064_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1186_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1594_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0063_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1187_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1595_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0061_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1188_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1596_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0062_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1189_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1597_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1186_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1187_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1188_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1189_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1190_ ) );
NOR2_X4 \u1_ps2_dsh/key_ascii/i0/_1598_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1185_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1190_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1191_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1599_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0295_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1192_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1600_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0294_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1193_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1601_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0290_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1194_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1602_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0289_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1195_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1603_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1192_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1193_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1194_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1195_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1196_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1604_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0291_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1197_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1605_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0287_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1198_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1606_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0292_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1199_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1607_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0288_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1200_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1608_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1197_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1198_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1199_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1200_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1201_ ) );
NOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1609_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1196_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1201_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1202_ ) );
NOR4_X1 \u1_ps2_dsh/key_ascii/i0/_1610_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1169_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1180_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1203_ ) );
NAND4_X2 \u1_ps2_dsh/key_ascii/i0/_1611_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1027_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1115_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1158_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1203_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1204_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1612_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0366_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1205_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1613_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0365_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1206_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1614_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0362_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1207_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1615_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0361_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1208_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1616_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1205_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1206_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1207_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1208_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1209_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1617_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0363_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1210_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1618_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0358_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1211_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1619_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0364_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1212_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1620_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0359_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1213_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1621_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1210_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1211_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1212_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1213_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1214_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1622_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1209_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1214_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1215_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1623_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0330_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1216_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1624_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0329_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1217_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1625_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0325_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1218_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1626_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0324_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1219_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1627_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1216_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1217_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1218_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1219_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1220_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1628_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0327_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1221_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1629_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0322_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1222_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1630_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0328_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1223_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1631_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0323_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1224_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1632_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1221_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1222_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1223_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1224_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1225_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1633_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1220_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1225_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1226_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1634_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0521_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1227_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1635_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0520_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1228_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1636_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0525_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1229_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1637_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0524_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1230_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1638_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1227_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1228_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1229_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1230_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1231_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1639_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0518_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1232_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1640_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0522_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1233_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1641_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0519_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1234_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1642_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0523_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1235_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1643_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1232_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1233_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1234_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1235_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1236_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1644_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1237_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1645_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0401_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1238_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1646_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0400_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1239_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1647_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0397_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1240_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1648_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0396_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1241_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1649_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1238_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1239_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1240_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1241_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1242_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1650_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0398_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1243_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1651_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0394_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1244_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1652_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0399_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1245_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1653_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0395_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1246_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1654_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1243_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1244_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1245_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1246_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1247_ ) );
NOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1655_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1242_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1247_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1248_ ) );
NOR4_X1 \u1_ps2_dsh/key_ascii/i0/_1656_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1215_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1226_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1237_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1249_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1657_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0436_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1250_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1658_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0435_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1251_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1659_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0433_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1252_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1660_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0434_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1253_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1661_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1250_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1251_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1252_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1253_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1254_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1662_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0432_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1255_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1663_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0431_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1256_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1664_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0429_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1257_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1665_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0430_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1258_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1666_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1255_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1256_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1257_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1258_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1259_ ) );
NOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1667_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1254_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1259_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1260_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1668_ ( .A(fanout_net_27 ), .B(\u1_ps2_dsh/key_ascii/i0/_0260_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1261_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1669_ ( .A(fanout_net_26 ), .B(\u1_ps2_dsh/key_ascii/i0/_0249_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1262_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1670_ ( .A(fanout_net_23 ), .B(\u1_ps2_dsh/key_ascii/i0/_0215_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1263_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1671_ ( .A(fanout_net_22 ), .B(\u1_ps2_dsh/key_ascii/i0/_0204_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1264_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1672_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1261_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1262_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1263_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1264_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1265_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1673_ ( .A(fanout_net_24 ), .B(\u1_ps2_dsh/key_ascii/i0/_0226_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1266_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1674_ ( .A(fanout_net_20 ), .B(\u1_ps2_dsh/key_ascii/i0/_0182_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1267_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1675_ ( .A(fanout_net_25 ), .B(\u1_ps2_dsh/key_ascii/i0/_0237_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1268_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1676_ ( .A(fanout_net_21 ), .B(\u1_ps2_dsh/key_ascii/i0/_0193_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1269_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1677_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1266_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1267_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1268_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1269_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1270_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1678_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1271_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1679_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0308_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1272_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1680_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0307_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1273_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1681_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0312_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1274_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1682_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0311_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1275_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1683_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1272_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1273_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1274_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1275_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1276_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1684_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0305_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1277_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1685_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0309_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1278_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1686_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0306_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1279_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1687_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0310_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1280_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1688_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1277_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1278_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1279_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1280_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1281_ ) );
AND2_X2 \u1_ps2_dsh/key_ascii/i0/_1689_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1276_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1281_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1282_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1690_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0586_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1283_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1691_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0585_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1284_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1692_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0582_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1285_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1693_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0581_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1286_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1694_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1283_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1284_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1285_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1286_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1287_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1695_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0583_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1288_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1696_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0578_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1289_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1697_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0584_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1290_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1698_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0579_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1291_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1699_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1288_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1289_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1290_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1291_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1292_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1700_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1293_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1701_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0343_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1294_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1702_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0342_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1295_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1703_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0347_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1296_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1704_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0346_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1297_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1705_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1294_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1295_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1296_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1297_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1298_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1706_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0340_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1299_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1707_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0344_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1300_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1708_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0341_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1301_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1709_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0345_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1302_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1710_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1299_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1300_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1301_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1302_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1303_ ) );
NOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1711_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1298_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1303_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1304_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1712_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0273_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1305_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1713_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0272_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1306_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1714_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0269_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1307_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1715_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0270_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1308_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1716_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1305_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1306_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1307_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1308_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1309_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1717_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0277_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1310_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1718_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0276_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1311_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1719_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0274_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1312_ ) );
XNOR2_X2 \u1_ps2_dsh/key_ascii/i0/_1720_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0275_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1313_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1721_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1310_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1311_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1312_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1313_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1314_ ) );
NOR2_X4 \u1_ps2_dsh/key_ascii/i0/_1722_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1309_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1314_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1315_ ) );
NOR4_X1 \u1_ps2_dsh/key_ascii/i0/_1723_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1293_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1316_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1724_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0117_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1317_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1725_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0116_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1318_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1726_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0112_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1319_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1727_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0111_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1320_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1728_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1317_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1318_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1319_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1320_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1321_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1729_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0113_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1322_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1730_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0109_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1323_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1731_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0114_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1324_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1732_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0110_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1325_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1733_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1322_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1323_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1324_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1325_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1326_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1734_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0082_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1327_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1735_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0071_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1328_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1736_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0038_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1329_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1737_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0027_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1330_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1738_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1327_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1328_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1329_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1330_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1331_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1739_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0049_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1332_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1740_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0580_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1333_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1741_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0060_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1334_ ) );
XNOR2_X1 \u1_ps2_dsh/key_ascii/i0/_1742_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .B(\u1_ps2_dsh/key_ascii/i0/_0591_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1335_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1743_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1332_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1333_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1334_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_1335_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0592_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1744_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0593_ ) );
NAND4_X4 \u1_ps2_dsh/key_ascii/i0/_1745_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1249_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1271_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_1316_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0593_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0594_ ) );
NOR2_X4 \u1_ps2_dsh/key_ascii/i0/_1746_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1204_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0594_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0595_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1747_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0000_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0596_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1748_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0509_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0597_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1749_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0438_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0598_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1750_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0598_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0992_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0402_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0474_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0969_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0599_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1751_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0296_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0261_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0600_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1752_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0367_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0601_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1753_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0597_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0599_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0600_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0601_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0602_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1754_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0278_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0603_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1755_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0385_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0604_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1756_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1220_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1225_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0313_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0605_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1757_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1209_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1214_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0350_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0606_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1758_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0603_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0604_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0605_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0606_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0607_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1759_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0243_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0608_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1760_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0030_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0609_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1761_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0570_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0610_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1762_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0207_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0611_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1763_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0608_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0609_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0610_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0611_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0612_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1764_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0587_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0613_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1765_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0552_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0614_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1766_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0271_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0615_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1767_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0016_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0616_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1768_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0613_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0614_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0615_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0616_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0617_ ) );
NOR3_X1 \u1_ps2_dsh/key_ascii/i0/_1769_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0607_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0612_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0617_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0618_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1770_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0224_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0619_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1771_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0189_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0620_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1772_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0118_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0621_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1773_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0154_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0622_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1774_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0619_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0620_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0621_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0622_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0623_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1775_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0448_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0624_ ) );
AND3_X2 \u1_ps2_dsh/key_ascii/i0/_1776_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0093_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0625_ ) );
OR2_X1 \u1_ps2_dsh/key_ascii/i0/_1777_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0624_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0625_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0626_ ) );
AOI221_X1 \u1_ps2_dsh/key_ascii/i0/_1778_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0626_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0047_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0083_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_1180_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0627_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1779_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0491_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0628_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1780_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0527_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0629_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1781_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0628_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0629_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0630_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1782_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0631_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1783_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0630_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0420_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0455_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0631_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0632_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1784_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0136_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0633_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1785_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0065_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0634_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1786_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0172_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0635_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1787_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0100_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0636_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1788_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0633_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0634_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0635_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0636_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0637_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_1789_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0623_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0627_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0632_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0637_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0638_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1790_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0596_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0602_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0618_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0638_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1336_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1791_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0001_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0639_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1792_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0510_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0640_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1793_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0475_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0641_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1794_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0641_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0992_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0403_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0439_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0947_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0642_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1795_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0297_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0262_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0643_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1796_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0332_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0368_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0644_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1797_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0640_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0642_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0643_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0644_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0645_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1798_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1220_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1225_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0314_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0646_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1799_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0646_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0279_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0647_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1800_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0244_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0648_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1801_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0208_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0649_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1802_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0031_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0650_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1803_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0571_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0651_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1804_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0648_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0649_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0650_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0651_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0652_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1805_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0282_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0653_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1806_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0127_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0654_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1807_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0553_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0655_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1808_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0588_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0656_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1809_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0653_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0654_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0655_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0656_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0657_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1810_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1215_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0351_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0386_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0658_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1811_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0647_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0652_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0657_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0658_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0659_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1812_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0155_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0660_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1813_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0119_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0661_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1814_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0190_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0662_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1815_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0225_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0663_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1816_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0660_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0661_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0662_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0663_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0664_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1817_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0492_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0665_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1818_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0528_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0666_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1819_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0665_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0666_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0667_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1820_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0667_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0421_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0456_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0631_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0668_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1821_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0048_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0669_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1822_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0084_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0670_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1823_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0669_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0670_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0671_ ) );
AND2_X2 \u1_ps2_dsh/key_ascii/i0/_1824_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0672_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1825_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0671_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0104_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0672_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0459_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0958_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0673_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1826_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0137_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0674_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1827_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0066_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0675_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1828_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0173_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0676_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1829_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0101_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0677_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1830_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0674_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0675_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0676_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0677_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0678_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1831_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0664_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0668_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0673_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0678_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0679_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1832_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0639_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0645_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0659_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0679_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1337_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1833_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0002_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0680_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1834_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0529_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0681_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1835_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0494_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0682_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1836_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0139_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0683_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1837_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0440_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0684_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1838_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0681_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0682_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0683_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0684_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0685_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1839_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0422_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0686_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1840_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0280_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0687_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1841_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0032_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0688_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1842_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0572_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0689_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1843_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0686_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0687_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0688_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0689_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0690_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1844_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0511_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0691_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1845_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0476_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0692_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1846_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0691_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0692_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0693_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1847_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0263_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0333_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0694_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1848_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0685_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0690_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0693_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0694_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0695_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1849_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0050_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0696_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1850_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0696_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0085_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1180_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0697_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1851_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0672_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0115_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0387_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0698_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1852_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1209_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1214_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0352_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0699_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1853_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0067_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0700_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1854_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0699_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0700_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0701_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1855_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0701_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0298_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0316_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_1226_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0702_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1856_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0697_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0698_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0702_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0703_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1857_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0369_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0704_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1858_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0120_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0705_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1859_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0457_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0706_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1860_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0245_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0707_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1861_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0704_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0705_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0706_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0707_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0708_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1862_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0209_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0709_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1863_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0238_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0710_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1864_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0554_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0711_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1865_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0293_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0712_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1866_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0709_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0710_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0711_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0712_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0713_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1867_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0227_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0714_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1868_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0471_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0715_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1869_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0191_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0716_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1870_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0156_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0717_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1871_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0714_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0715_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0716_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0717_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0718_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1872_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0174_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0719_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1873_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0589_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0720_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1874_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0986_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0991_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0405_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0721_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1875_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0102_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0722_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1876_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0719_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0720_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0721_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0722_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0723_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1877_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0708_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0713_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0718_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0723_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0724_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1878_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0680_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0695_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0703_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0724_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1338_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1879_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0003_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0725_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1880_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0192_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0726_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1881_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0512_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0727_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1882_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0441_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0728_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1883_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0477_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0729_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1884_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0986_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0991_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0406_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0730_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1885_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0727_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0728_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0729_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0730_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0731_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1886_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0121_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0732_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1887_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0157_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0733_ ) );
AND2_X1 \u1_ps2_dsh/key_ascii/i0/_1888_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0732_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0733_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0734_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1889_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0980_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0228_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0370_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0735_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1890_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0726_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0731_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0734_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0735_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0736_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1891_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1215_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0353_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0388_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0737_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1892_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0210_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0738_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1893_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0573_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0739_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1894_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0246_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0740_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1895_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0033_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0741_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1896_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0738_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0739_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0740_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0741_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0742_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1897_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0349_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0743_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1898_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0590_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0744_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1899_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0555_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0745_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1900_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0304_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0746_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1901_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0743_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0744_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0745_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0746_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0747_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1902_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1226_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0317_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0281_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0748_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1903_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0737_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0742_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0747_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0748_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0749_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1904_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1276_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1281_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0299_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0750_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1905_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0750_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0264_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0334_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0751_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1906_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0051_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0752_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1907_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0086_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0753_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1908_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0752_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0753_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0754_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_1909_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0754_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0126_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0672_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0482_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0958_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0755_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1910_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0423_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0756_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1911_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0495_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0757_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1912_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0530_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0758_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1913_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0458_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0759_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1914_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0756_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0757_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0758_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0759_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0760_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1915_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0103_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0761_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1916_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0140_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0762_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1917_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0068_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0763_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1918_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0175_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0764_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1919_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0761_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0762_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0763_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0764_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0765_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_1920_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0751_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0755_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0760_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0765_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0766_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1921_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0725_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0736_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0749_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0766_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1339_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1922_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0004_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0767_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1923_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0513_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0768_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1924_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0986_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0991_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0407_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0769_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1925_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0478_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0770_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1926_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0442_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0771_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1927_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0768_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0769_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0770_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0771_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0772_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1928_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0300_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0265_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0773_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1929_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0335_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0372_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0774_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1930_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0772_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0773_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0774_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0775_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1931_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0496_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0776_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1932_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0461_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0777_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1933_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0531_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0778_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1934_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0776_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0777_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0778_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0779_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1935_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0460_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0780_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1936_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0017_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0781_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1937_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0556_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0782_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1938_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0783_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1939_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0780_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0781_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0782_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0783_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0784_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1940_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0283_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0424_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0785_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1941_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0211_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0786_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1942_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0574_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0787_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1943_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0247_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0788_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1944_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0034_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0789_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1945_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0786_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0787_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0788_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0789_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0790_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1946_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0779_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0784_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0785_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0790_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0791_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1947_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0141_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0792_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1948_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0105_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0793_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1949_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0069_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0794_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1950_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0176_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0795_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1951_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0792_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0793_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0794_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0795_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0796_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1952_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0052_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0797_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1953_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0493_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0798_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1954_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0087_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0799_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1955_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0138_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0800_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1956_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0797_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0798_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0799_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0800_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0801_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1957_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0158_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0802_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1958_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0122_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0803_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1959_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0194_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0804_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1960_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0229_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0805_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1961_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0802_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0803_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0804_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0805_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0806_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1962_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0389_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0807_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1963_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1220_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1225_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0318_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0808_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1964_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1209_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1214_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0354_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0809_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1965_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0807_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0808_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0809_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0810_ ) );
NOR4_X1 \u1_ps2_dsh/key_ascii/i0/_1966_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0796_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0801_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0806_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0810_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0811_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_1967_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0767_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0775_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0791_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0811_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1340_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1968_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0005_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0812_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_1969_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0159_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0813_ ) );
AOI21_X1 \u1_ps2_dsh/key_ascii/i0/_1970_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0813_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0123_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1003_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0814_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1971_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0479_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0815_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1972_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0514_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0816_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1973_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0941_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0946_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0443_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0817_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1974_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0986_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0991_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0408_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0818_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1975_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0815_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0816_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0817_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0818_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0819_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1976_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0195_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0820_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1977_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0980_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0230_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0373_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0821_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1978_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0814_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0819_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0820_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0821_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0822_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1979_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1215_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0355_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0390_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0823_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1980_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0824_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1981_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0575_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0825_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1982_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0212_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0826_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1983_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0035_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0827_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1984_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0824_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0825_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0826_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0827_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0828_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1985_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0547_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0829_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1986_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0557_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0830_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1987_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0326_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0831_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1988_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0018_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0832_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1989_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0829_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0830_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0831_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0832_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0833_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_1990_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1226_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0319_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0284_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0834_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1991_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0823_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0828_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0833_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0834_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0835_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1992_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0106_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0836_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1993_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0142_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0837_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1994_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0070_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0838_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1995_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0177_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0839_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_1996_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0836_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0837_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0838_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0839_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0840_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1997_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0149_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0841_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_1998_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0504_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0842_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_1999_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0841_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0842_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0843_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_2000_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0843_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0053_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0088_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_1180_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0844_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2001_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0425_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0845_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2002_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0497_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0846_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2003_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0462_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0847_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2004_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0532_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0848_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2005_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0845_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0846_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0847_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0848_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0849_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_2006_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1276_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1281_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0301_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0850_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_2007_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0850_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0266_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0336_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0851_ ) );
AND4_X2 \u1_ps2_dsh/key_ascii/i0/_2008_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0840_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0844_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0849_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0851_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0852_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2009_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0812_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0822_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0835_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0852_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1341_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2010_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0006_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0853_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2011_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0516_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0854_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_2012_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0480_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0855_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_2013_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0855_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0992_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0409_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0444_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0947_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0856_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2014_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0302_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0267_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0857_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2015_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0338_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0374_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0858_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2016_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0854_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0856_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0857_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0858_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0859_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2017_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1215_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0356_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0391_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0860_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2018_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0250_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0861_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2019_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0036_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0862_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2020_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0213_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0863_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2021_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0576_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0864_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2022_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0861_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0862_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0863_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0864_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0865_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2023_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0558_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0866_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2024_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0337_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0867_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2025_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0559_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0868_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2026_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0019_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0869_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2027_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0866_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0867_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0868_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0869_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0870_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2028_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1226_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0320_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0285_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0871_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2029_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0860_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0865_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0870_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0871_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0872_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2030_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0161_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0873_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2031_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0124_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0874_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2032_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0196_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0875_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2033_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0231_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0876_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2034_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0873_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0874_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0875_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0876_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0877_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2035_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0089_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0878_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2036_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0054_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0879_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2037_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0952_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0957_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0515_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0880_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2038_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1265_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1270_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0160_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0881_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2039_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0878_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0879_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0880_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0881_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0882_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2040_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0427_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0883_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2041_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0498_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0884_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2042_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0533_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0885_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2043_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0463_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0886_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2044_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0883_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0884_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0885_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0886_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0887_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2045_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0107_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0888_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2046_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0143_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0889_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2047_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0072_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0890_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2048_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0178_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0891_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2049_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0888_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0889_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0890_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0891_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0892_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2050_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0877_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0882_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0887_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0892_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0893_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2051_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0853_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0859_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0872_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0893_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1342_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2052_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0595_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0007_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0894_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2053_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1231_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1236_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0517_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0895_ ) );
AND3_X1 \u1_ps2_dsh/key_ascii/i0/_2054_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0963_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0968_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0481_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0896_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_2055_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0896_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0992_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0410_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0445_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0947_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0897_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2056_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1282_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0303_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0268_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_1315_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0898_ ) );
AOI22_X1 \u1_ps2_dsh/key_ascii/i0/_2057_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0339_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1304_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_1015_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0375_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0899_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2058_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0895_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0897_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0898_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0899_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0900_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2059_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1202_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0286_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0901_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2060_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1248_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0392_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0902_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2061_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1220_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1225_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0321_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0903_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2062_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1209_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1214_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0357_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0904_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2063_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0901_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0902_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0903_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0904_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0905_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2064_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1064_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1069_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0251_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0906_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2065_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1141_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1146_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0037_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0907_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2066_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1287_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1292_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0577_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0908_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2067_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1032_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1037_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0214_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0909_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2068_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0906_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0907_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0908_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0909_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0910_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2069_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1163_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1168_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0020_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0911_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2070_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1130_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1135_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0560_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0912_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2071_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1151_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1156_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0348_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0913_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2072_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1331_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0592_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0569_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0914_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2073_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0911_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0912_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0913_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0914_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0915_ ) );
NOR3_X1 \u1_ps2_dsh/key_ascii/i0/_2074_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0905_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0910_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0915_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0916_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2075_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0974_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0979_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0232_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0917_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2076_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1086_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1091_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0197_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0918_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2077_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0997_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1002_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0125_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0919_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2078_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1020_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1025_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0162_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0920_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2079_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0917_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0918_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0919_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0920_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0921_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2080_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1191_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0055_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0922_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2081_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1174_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1179_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0090_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0923_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2082_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0922_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0923_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0924_ ) );
AOI221_X4 \u1_ps2_dsh/key_ascii/i0/_2083_ ( .A(\u1_ps2_dsh/key_ascii/i0/_0924_ ), .B1(\u1_ps2_dsh/key_ascii/i0/_0171_ ), .B2(\u1_ps2_dsh/key_ascii/i0/_0672_ ), .C1(\u1_ps2_dsh/key_ascii/i0/_0526_ ), .C2(\u1_ps2_dsh/key_ascii/i0/_0958_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0925_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2084_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1081_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0499_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0926_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2085_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1260_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0428_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0927_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2086_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1054_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1059_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0464_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0928_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2087_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1108_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1113_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0534_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0929_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2088_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0926_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0927_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0928_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0929_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0930_ ) );
NAND2_X1 \u1_ps2_dsh/key_ascii/i0/_2089_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1103_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0144_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0931_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2090_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1321_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1326_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0108_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0932_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2091_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1043_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1048_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0179_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0933_ ) );
NAND3_X1 \u1_ps2_dsh/key_ascii/i0/_2092_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_1120_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_1125_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0073_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0934_ ) );
AND4_X1 \u1_ps2_dsh/key_ascii/i0/_2093_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0931_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0932_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0933_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0934_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0935_ ) );
AND4_X4 \u1_ps2_dsh/key_ascii/i0/_2094_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0921_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0925_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0930_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0935_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_0936_ ) );
NAND4_X1 \u1_ps2_dsh/key_ascii/i0/_2095_ ( .A1(\u1_ps2_dsh/key_ascii/i0/_0894_ ), .A2(\u1_ps2_dsh/key_ascii/i0/_0900_ ), .A3(\u1_ps2_dsh/key_ascii/i0/_0916_ ), .A4(\u1_ps2_dsh/key_ascii/i0/_0936_ ), .ZN(\u1_ps2_dsh/key_ascii/i0/_1343_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2096_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0535_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2097_ ( .A(\data_d1 [0] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0008_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2098_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0536_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2099_ ( .A(\data_d1 [1] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0009_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2100_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0538_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2101_ ( .A(\data_d1 [2] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0010_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2102_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0539_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2103_ ( .A(\data_d1 [3] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0011_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2104_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0540_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2105_ ( .A(\data_d1 [4] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0012_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2106_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0541_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2107_ ( .A(\data_d1 [5] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0013_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2108_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0542_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2109_ ( .A(\data_d1 [6] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0014_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2110_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0543_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2111_ ( .A(\data_d1 [7] ), .Z(\u1_ps2_dsh/key_ascii/i0/_0015_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2112_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0518_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2113_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0519_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2114_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0520_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2115_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0521_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2116_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0522_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2117_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0523_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2118_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0524_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2119_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0525_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2120_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0500_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2121_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0501_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2122_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0502_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2123_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0503_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2124_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0505_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2125_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0506_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2126_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0507_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2127_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0508_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2128_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0483_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2129_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0484_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2130_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0485_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2131_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0486_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2132_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0487_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2133_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0488_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2134_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0489_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2135_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0490_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2136_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0465_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2137_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0466_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2138_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0467_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2139_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0468_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2140_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0469_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2141_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0470_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2142_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0472_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2143_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0473_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2144_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0446_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2145_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0447_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2146_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0449_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2147_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0450_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2148_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0451_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2149_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0452_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2150_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0453_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2151_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0454_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2152_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0429_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2153_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0430_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2154_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0431_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2155_ ( .A(fanout_net_9 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0432_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2156_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0433_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2157_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0434_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2158_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0435_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2159_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0436_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2160_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0411_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2161_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0412_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2162_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0413_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2163_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0414_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2164_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0416_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2165_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0417_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2166_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0418_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2167_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0419_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2168_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0394_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2169_ ( .A(fanout_net_1 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0395_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2170_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0396_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2171_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0397_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2172_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0398_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2173_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0399_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2174_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0400_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2175_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0401_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2176_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0376_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2177_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0377_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2178_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0378_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2179_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0379_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2180_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0380_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2181_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0381_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2182_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0383_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2183_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0384_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2184_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0358_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2185_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0359_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2186_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0361_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2187_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0362_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2188_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0363_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2189_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0364_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2190_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0365_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2191_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0366_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2192_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0340_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2193_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0341_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2194_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0342_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2195_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0343_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2196_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0344_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2197_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0345_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2198_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0346_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2199_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0347_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2200_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0322_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2201_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0323_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2202_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0324_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2203_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0325_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2204_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0327_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2205_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0328_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2206_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0329_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2207_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0330_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2208_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0305_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2209_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0306_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2210_ ( .A(fanout_net_10 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0307_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2211_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0308_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2212_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0309_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2213_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0310_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2214_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0311_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2215_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0312_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2216_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0287_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2217_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0288_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2218_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0289_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2219_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0290_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2220_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0291_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2221_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0292_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2222_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0294_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2223_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0295_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2224_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0269_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2225_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0270_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2226_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0272_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2227_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0273_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2228_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0274_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2229_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0275_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2230_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0276_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2231_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0277_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2232_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0252_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2233_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0253_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2234_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0254_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2235_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0255_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2236_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0256_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2237_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0257_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2238_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0258_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2239_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0259_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2240_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0233_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2241_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0234_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2242_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0235_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2243_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0236_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2244_ ( .A(fanout_net_2 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0239_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2245_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0240_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2246_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0241_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2247_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0242_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2248_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0216_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2249_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0217_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2250_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0218_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2251_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0219_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2252_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0220_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2253_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0221_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2254_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0222_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2255_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0223_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2256_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0198_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2257_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0199_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2258_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0200_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2259_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0201_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2260_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0202_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2261_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0203_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2262_ ( .A(fanout_net_11 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0205_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2263_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0206_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2264_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0180_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2265_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0181_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2266_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0183_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2267_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0184_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2268_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0185_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2269_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0186_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2270_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0187_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2271_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0188_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2272_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0163_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2273_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0164_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2274_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0165_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2275_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0166_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2276_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0167_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2277_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0168_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2278_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0169_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2279_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0170_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2280_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0145_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2281_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0146_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2282_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0147_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2283_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0148_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2284_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0150_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2285_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0151_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2286_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0152_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2287_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0153_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2288_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0128_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2289_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0129_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2290_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0130_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2291_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0131_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2292_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0132_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2293_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0133_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2294_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0134_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2295_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0135_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2296_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0109_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2297_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0110_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2298_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0111_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2299_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0112_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2300_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0113_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2301_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0114_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2302_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0116_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2303_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0117_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2304_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0091_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2305_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0092_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2306_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0094_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2307_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0095_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2308_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0096_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2309_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0097_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2310_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0098_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2311_ ( .A(fanout_net_12 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0099_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2312_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0074_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2313_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0075_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2314_ ( .A(fanout_net_3 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0076_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2315_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0077_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2316_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0078_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2317_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0079_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2318_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0080_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2319_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0081_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2320_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0056_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2321_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0057_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2322_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0058_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2323_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0059_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2324_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0061_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2325_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0062_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2326_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0063_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2327_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0064_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2328_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0039_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2329_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0040_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2330_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0041_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2331_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0042_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2332_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0043_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2333_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0044_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2334_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0045_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2335_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0046_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2336_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0021_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2337_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0022_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2338_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0023_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2339_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0024_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2340_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0025_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2341_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0026_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2342_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0028_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2343_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0029_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2344_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0578_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2345_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0579_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2346_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0581_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2347_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0582_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2348_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0583_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2349_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0584_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2350_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0585_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2351_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0586_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2352_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0561_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2353_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0562_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2354_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0563_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2355_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0564_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2356_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0565_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2357_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0566_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2358_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0567_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2359_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0568_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2360_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0537_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2361_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0544_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2362_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0545_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2363_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0546_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2364_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0548_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2365_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0549_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2366_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0550_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2367_ ( .A(fanout_net_13 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0551_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2368_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0360_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2369_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0371_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2370_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0382_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2371_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0393_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2372_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0404_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2373_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0415_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2374_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0426_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2375_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0437_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2376_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0580_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2377_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0591_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2378_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0027_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2379_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0038_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2380_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0049_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2381_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0060_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2382_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0071_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2383_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0082_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2384_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0182_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2385_ ( .A(fanout_net_4 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0193_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2386_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0204_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2387_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0215_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2388_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0226_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2389_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0237_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2390_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0249_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2391_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0260_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2392_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0016_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2393_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0093_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2394_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0271_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2395_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0448_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2396_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0552_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2397_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0570_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2398_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0587_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2399_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0030_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2400_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0047_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2401_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0065_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2402_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0083_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2403_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0100_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2404_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0118_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2405_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0136_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2406_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0154_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2407_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0172_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2408_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0189_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2409_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0207_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2410_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0224_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2411_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0243_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2412_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0261_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2413_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0278_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2414_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0296_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2415_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0313_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2416_ ( .A(fanout_net_14 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0331_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2417_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0350_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2418_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0367_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2419_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0385_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2420_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0402_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2421_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0420_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2422_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0438_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2423_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0455_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2424_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0474_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2425_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0491_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2426_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0509_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2427_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0527_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2428_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0000_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2429_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1336_ ), .Z(\u1_ps2_dsh/ascii_result [0] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2430_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0127_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2431_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0104_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2432_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0282_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2433_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0459_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2434_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0553_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2435_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0571_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2436_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0588_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2437_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0031_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2438_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0048_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2439_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0066_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2440_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0084_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2441_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0101_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2442_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0119_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2443_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0137_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2444_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0155_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2445_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0173_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2446_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0190_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2447_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0208_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2448_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0225_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2449_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0244_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2450_ ( .A(fanout_net_5 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0262_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2451_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0279_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2452_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0297_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2453_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0314_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2454_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0332_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2455_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0351_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2456_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0368_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2457_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0386_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2458_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0403_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2459_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0421_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2460_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0439_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2461_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0456_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2462_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0475_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2463_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0492_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2464_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0510_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2465_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0528_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2466_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0001_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2467_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1337_ ), .Z(\u1_ps2_dsh/ascii_result [1] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2468_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0238_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2469_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0115_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2470_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0293_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2471_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0471_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2472_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0554_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2473_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0572_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2474_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0589_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2475_ ( .A(fanout_net_15 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0032_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2476_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0050_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2477_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0067_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2478_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0085_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2479_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0102_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2480_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0120_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2481_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0139_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2482_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0156_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2483_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0174_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2484_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0191_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2485_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0209_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2486_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0227_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2487_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0245_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2488_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0263_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2489_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0280_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2490_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0298_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2491_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0316_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2492_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0333_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2493_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0352_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2494_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0369_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2495_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0387_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2496_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0405_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2497_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0422_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2498_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0440_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2499_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0457_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2500_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0476_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2501_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0494_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2502_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0511_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2503_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0529_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2504_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0002_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2505_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1338_ ), .Z(\u1_ps2_dsh/ascii_result [2] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2506_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0349_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2507_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0126_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2508_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0304_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2509_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0482_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2510_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0555_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2511_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0573_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2512_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0590_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2513_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0033_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2514_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0051_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2515_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0068_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2516_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0086_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2517_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0103_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2518_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0121_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2519_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0140_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2520_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0157_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2521_ ( .A(fanout_net_6 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0175_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2522_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0192_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2523_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0210_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2524_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0228_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2525_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0246_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2526_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0264_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2527_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0281_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2528_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0299_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2529_ ( .A(fanout_net_16 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0317_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2530_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0334_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2531_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0353_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2532_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0370_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2533_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0388_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2534_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0406_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2535_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0423_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2536_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0441_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2537_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0458_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2538_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0477_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2539_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0495_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2540_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0512_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2541_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0530_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2542_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0003_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2543_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1339_ ), .Z(\u1_ps2_dsh/ascii_result [3] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2544_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0460_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2545_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0138_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2546_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0315_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2547_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0493_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2548_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0556_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2549_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0574_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2550_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0017_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2551_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0034_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2552_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0052_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2553_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0069_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2554_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0087_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2555_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0105_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2556_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0122_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2557_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0141_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2558_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0158_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2559_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0176_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2560_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0194_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2561_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0211_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2562_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0229_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2563_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0247_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2564_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0265_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2565_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0283_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2566_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0300_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2567_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0318_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2568_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0335_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2569_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0354_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2570_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0372_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2571_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0389_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2572_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0407_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2573_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0424_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2574_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0442_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2575_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0461_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2576_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0478_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2577_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0496_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2578_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0513_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2579_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0531_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2580_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0004_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2581_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1340_ ), .Z(\u1_ps2_dsh/ascii_result [4] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2582_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0547_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2583_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0149_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2584_ ( .A(fanout_net_17 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0326_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2585_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0504_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2586_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0557_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2587_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0575_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2588_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0018_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2589_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0035_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2590_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0053_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2591_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0070_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2592_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0088_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2593_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0106_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2594_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0123_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2595_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0142_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2596_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0159_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2597_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0177_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2598_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0195_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2599_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0212_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2600_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0230_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2601_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0248_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2602_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0266_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2603_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0284_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2604_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0301_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2605_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0319_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2606_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0336_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2607_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0355_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2608_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0373_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2609_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0390_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2610_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0408_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2611_ ( .A(fanout_net_7 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0425_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2612_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0443_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2613_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0462_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2614_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0479_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2615_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0497_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2616_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0514_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2617_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0532_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2618_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0005_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2619_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1341_ ), .Z(\u1_ps2_dsh/ascii_result [5] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2620_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0558_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2621_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0160_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2622_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0337_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2623_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0515_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2624_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0559_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2625_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0576_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2626_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0019_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2627_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0036_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2628_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0054_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2629_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0072_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2630_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0089_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2631_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0107_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2632_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0124_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2633_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0143_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2634_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0161_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2635_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0178_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2636_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0196_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2637_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0213_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2638_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0231_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2639_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0250_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2640_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0267_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2641_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0285_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2642_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0302_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2643_ ( .A(fanout_net_8 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0320_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2644_ ( .A(\u1_ps2_dsh/_050_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0338_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2645_ ( .A(\u1_ps2_dsh/_050_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0356_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2646_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0374_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2647_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0391_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2648_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0409_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2649_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0427_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2650_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0444_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2651_ ( .A(fanout_net_18 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0463_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2652_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0480_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2653_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0498_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2654_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0516_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2655_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0533_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2656_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0006_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2657_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1342_ ), .Z(\u1_ps2_dsh/ascii_result [6] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2658_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0569_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2659_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0171_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2660_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0348_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2661_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0526_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2662_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0560_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2663_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0577_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2664_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0020_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2665_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0037_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2666_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0055_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2667_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0073_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2668_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0090_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2669_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0108_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2670_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0125_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2671_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0144_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2672_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0162_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2673_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0179_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2674_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0197_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2675_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0214_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2676_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0232_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2677_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0251_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2678_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0268_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2679_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0286_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2680_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0303_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2681_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0321_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2682_ ( .A(fanout_net_19 ), .Z(\u1_ps2_dsh/key_ascii/i0/_0339_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2683_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0357_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2684_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0375_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2685_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0392_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2686_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0410_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2687_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0428_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2688_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0445_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2689_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0464_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2690_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0481_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2691_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0499_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2692_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0517_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2693_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0534_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2694_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/key_ascii/i0/_0007_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2695_ ( .A(\u1_ps2_dsh/key_ascii/i0/_1343_ ), .Z(\u1_ps2_dsh/ascii_result [7] ) );
INV_X32 \u2_ps2_cer/_067_ ( .A(\u2_ps2_cer/_056_ ), .ZN(\u2_ps2_cer/_021_ ) );
AND2_X4 \u2_ps2_cer/_068_ ( .A1(\u2_ps2_cer/_021_ ), .A2(\u2_ps2_cer/_057_ ), .ZN(\u2_ps2_cer/_022_ ) );
INV_X32 \u2_ps2_cer/_069_ ( .A(\u2_ps2_cer/_054_ ), .ZN(\u2_ps2_cer/_023_ ) );
NOR2_X4 \u2_ps2_cer/_070_ ( .A1(\u2_ps2_cer/_023_ ), .A2(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_024_ ) );
AND2_X4 \u2_ps2_cer/_071_ ( .A1(\u2_ps2_cer/_022_ ), .A2(\u2_ps2_cer/_024_ ), .ZN(\u2_ps2_cer/_025_ ) );
INV_X32 \u2_ps2_cer/_072_ ( .A(\u2_ps2_cer/_018_ ), .ZN(\u2_ps2_cer/_026_ ) );
AND2_X4 \u2_ps2_cer/_073_ ( .A1(\u2_ps2_cer/_026_ ), .A2(\u2_ps2_cer/_019_ ), .ZN(\u2_ps2_cer/_027_ ) );
AND2_X4 \u2_ps2_cer/_074_ ( .A1(\u2_ps2_cer/_025_ ), .A2(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_028_ ) );
INV_X16 \u2_ps2_cer/_075_ ( .A(\u2_ps2_cer/_050_ ), .ZN(\u2_ps2_cer/_029_ ) );
XNOR2_X1 \u2_ps2_cer/_076_ ( .A(\u2_ps2_cer/_028_ ), .B(\u2_ps2_cer/_029_ ), .ZN(\u2_ps2_cer/_010_ ) );
NOR2_X1 \u2_ps2_cer/_077_ ( .A1(\u2_ps2_cer/_029_ ), .A2(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_030_ ) );
INV_X2 \u2_ps2_cer/_078_ ( .A(\u2_ps2_cer/_053_ ), .ZN(\u2_ps2_cer/_031_ ) );
OAI211_X2 \u2_ps2_cer/_079_ ( .A(\u2_ps2_cer/_028_ ), .B(\u2_ps2_cer/_030_ ), .C1(\u2_ps2_cer/_052_ ), .C2(\u2_ps2_cer/_031_ ), .ZN(\u2_ps2_cer/_032_ ) );
INV_X1 \u2_ps2_cer/_080_ ( .A(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_033_ ) );
AND3_X1 \u2_ps2_cer/_081_ ( .A1(\u2_ps2_cer/_025_ ), .A2(\u2_ps2_cer/_050_ ), .A3(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_034_ ) );
OAI21_X1 \u2_ps2_cer/_082_ ( .A(\u2_ps2_cer/_032_ ), .B1(\u2_ps2_cer/_033_ ), .B2(\u2_ps2_cer/_034_ ), .ZN(\u2_ps2_cer/_011_ ) );
AND2_X4 \u2_ps2_cer/_083_ ( .A1(\u2_ps2_cer/_050_ ), .A2(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_035_ ) );
NAND2_X2 \u2_ps2_cer/_084_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_035_ ), .ZN(\u2_ps2_cer/_036_ ) );
XNOR2_X1 \u2_ps2_cer/_085_ ( .A(\u2_ps2_cer/_036_ ), .B(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_012_ ) );
NAND4_X1 \u2_ps2_cer/_086_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_052_ ), .A3(\u2_ps2_cer/_031_ ), .A4(\u2_ps2_cer/_035_ ), .ZN(\u2_ps2_cer/_037_ ) );
INV_X1 \u2_ps2_cer/_087_ ( .A(\u2_ps2_cer/_028_ ), .ZN(\u2_ps2_cer/_038_ ) );
NOR2_X1 \u2_ps2_cer/_088_ ( .A1(\u2_ps2_cer/_031_ ), .A2(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_039_ ) );
AOI22_X1 \u2_ps2_cer/_089_ ( .A1(\u2_ps2_cer/_039_ ), .A2(\u2_ps2_cer/_030_ ), .B1(\u2_ps2_cer/_035_ ), .B2(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_040_ ) );
NOR2_X2 \u2_ps2_cer/_090_ ( .A1(\u2_ps2_cer/_038_ ), .A2(\u2_ps2_cer/_040_ ), .ZN(\u2_ps2_cer/_041_ ) );
OAI21_X1 \u2_ps2_cer/_091_ ( .A(\u2_ps2_cer/_037_ ), .B1(\u2_ps2_cer/_041_ ), .B2(\u2_ps2_cer/_031_ ), .ZN(\u2_ps2_cer/_013_ ) );
XNOR2_X1 \u2_ps2_cer/_092_ ( .A(\u2_ps2_cer/_027_ ), .B(\u2_ps2_cer/_023_ ), .ZN(\u2_ps2_cer/_014_ ) );
NAND3_X1 \u2_ps2_cer/_093_ ( .A1(\u2_ps2_cer/_024_ ), .A2(\u2_ps2_cer/_026_ ), .A3(\u2_ps2_cer/_019_ ), .ZN(\u2_ps2_cer/_042_ ) );
AND3_X4 \u2_ps2_cer/_094_ ( .A1(\u2_ps2_cer/_026_ ), .A2(\u2_ps2_cer/_019_ ), .A3(\u2_ps2_cer/_054_ ), .ZN(\u2_ps2_cer/_043_ ) );
INV_X1 \u2_ps2_cer/_095_ ( .A(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_044_ ) );
OAI22_X1 \u2_ps2_cer/_096_ ( .A1(\u2_ps2_cer/_042_ ), .A2(\u2_ps2_cer/_022_ ), .B1(\u2_ps2_cer/_043_ ), .B2(\u2_ps2_cer/_044_ ), .ZN(\u2_ps2_cer/_015_ ) );
AND2_X4 \u2_ps2_cer/_097_ ( .A1(\u2_ps2_cer/_054_ ), .A2(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_045_ ) );
AND2_X2 \u2_ps2_cer/_098_ ( .A1(\u2_ps2_cer/_027_ ), .A2(\u2_ps2_cer/_045_ ), .ZN(\u2_ps2_cer/_046_ ) );
XNOR2_X1 \u2_ps2_cer/_099_ ( .A(\u2_ps2_cer/_046_ ), .B(\u2_ps2_cer/_021_ ), .ZN(\u2_ps2_cer/_016_ ) );
AOI21_X1 \u2_ps2_cer/_100_ ( .A(\u2_ps2_cer/_057_ ), .B1(\u2_ps2_cer/_046_ ), .B2(\u2_ps2_cer/_056_ ), .ZN(\u2_ps2_cer/_047_ ) );
AND4_X1 \u2_ps2_cer/_101_ ( .A1(\u2_ps2_cer/_056_ ), .A2(\u2_ps2_cer/_027_ ), .A3(\u2_ps2_cer/_057_ ), .A4(\u2_ps2_cer/_045_ ), .ZN(\u2_ps2_cer/_048_ ) );
NOR3_X1 \u2_ps2_cer/_102_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_047_ ), .A3(\u2_ps2_cer/_048_ ), .ZN(\u2_ps2_cer/_017_ ) );
INV_X1 \u2_ps2_cer/_103_ ( .A(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_049_ ) );
OAI21_X1 \u2_ps2_cer/_104_ ( .A(\u2_ps2_cer/_049_ ), .B1(\u2_ps2_cer/_026_ ), .B2(\u2_ps2_cer/_020_ ), .ZN(\u2_ps2_cer/_009_ ) );
BUF_X1 \u2_ps2_cer/_105_ ( .A(\u2_ps2_cer/counted ), .Z(\u2_ps2_cer/_018_ ) );
BUF_X1 \u2_ps2_cer/_106_ ( .A(_026_ ), .Z(\u2_ps2_cer/_019_ ) );
BUF_X1 \u2_ps2_cer/_107_ ( .A(\high_tens [0] ), .Z(\u2_ps2_cer/_050_ ) );
BUF_X1 \u2_ps2_cer/_108_ ( .A(\high_tens [1] ), .Z(\u2_ps2_cer/_051_ ) );
BUF_X1 \u2_ps2_cer/_109_ ( .A(\high_tens [2] ), .Z(\u2_ps2_cer/_052_ ) );
BUF_X1 \u2_ps2_cer/_110_ ( .A(\high_tens [3] ), .Z(\u2_ps2_cer/_053_ ) );
BUF_X1 \u2_ps2_cer/_111_ ( .A(\high_units [0] ), .Z(\u2_ps2_cer/_054_ ) );
BUF_X1 \u2_ps2_cer/_112_ ( .A(\high_units [1] ), .Z(\u2_ps2_cer/_055_ ) );
BUF_X1 \u2_ps2_cer/_113_ ( .A(\high_units [2] ), .Z(\u2_ps2_cer/_056_ ) );
BUF_X1 \u2_ps2_cer/_114_ ( .A(\high_units [3] ), .Z(\u2_ps2_cer/_057_ ) );
BUF_X1 \u2_ps2_cer/_115_ ( .A(\u2_ps2_cer/_010_ ), .Z(\u2_ps2_cer/_001_ ) );
BUF_X1 \u2_ps2_cer/_116_ ( .A(\u2_ps2_cer/_011_ ), .Z(\u2_ps2_cer/_002_ ) );
BUF_X1 \u2_ps2_cer/_117_ ( .A(\u2_ps2_cer/_012_ ), .Z(\u2_ps2_cer/_003_ ) );
BUF_X1 \u2_ps2_cer/_118_ ( .A(\u2_ps2_cer/_013_ ), .Z(\u2_ps2_cer/_004_ ) );
BUF_X1 \u2_ps2_cer/_119_ ( .A(\u2_ps2_cer/_014_ ), .Z(\u2_ps2_cer/_005_ ) );
BUF_X1 \u2_ps2_cer/_120_ ( .A(\u2_ps2_cer/_015_ ), .Z(\u2_ps2_cer/_006_ ) );
BUF_X1 \u2_ps2_cer/_121_ ( .A(\u2_ps2_cer/_016_ ), .Z(\u2_ps2_cer/_007_ ) );
BUF_X1 \u2_ps2_cer/_122_ ( .A(\u2_ps2_cer/_017_ ), .Z(\u2_ps2_cer/_008_ ) );
BUF_X1 \u2_ps2_cer/_123_ ( .A(key_release ), .Z(\u2_ps2_cer/_020_ ) );
BUF_X1 \u2_ps2_cer/_124_ ( .A(\u2_ps2_cer/_009_ ), .Z(\u2_ps2_cer/_000_ ) );
DFFR_X1 \u2_ps2_cer/_125_ ( .D(\u2_ps2_cer/_005_ ), .RN(clrn ), .CK(clk ), .Q(\high_units [0] ), .QN(\u2_ps2_cer/_058_ ) );
DFFR_X1 \u2_ps2_cer/_126_ ( .D(\u2_ps2_cer/_006_ ), .RN(clrn ), .CK(clk ), .Q(\high_units [1] ), .QN(\u2_ps2_cer/_059_ ) );
DFFR_X1 \u2_ps2_cer/_127_ ( .D(\u2_ps2_cer/_007_ ), .RN(clrn ), .CK(clk ), .Q(\high_units [2] ), .QN(\u2_ps2_cer/_060_ ) );
DFFR_X1 \u2_ps2_cer/_128_ ( .D(\u2_ps2_cer/_008_ ), .RN(clrn ), .CK(clk ), .Q(\high_units [3] ), .QN(\u2_ps2_cer/_061_ ) );
DFFR_X1 \u2_ps2_cer/_129_ ( .D(\u2_ps2_cer/_001_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens [0] ), .QN(\u2_ps2_cer/_062_ ) );
DFFR_X1 \u2_ps2_cer/_130_ ( .D(\u2_ps2_cer/_002_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens [1] ), .QN(\u2_ps2_cer/_063_ ) );
DFFR_X1 \u2_ps2_cer/_131_ ( .D(\u2_ps2_cer/_003_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens [2] ), .QN(\u2_ps2_cer/_064_ ) );
DFFR_X1 \u2_ps2_cer/_132_ ( .D(\u2_ps2_cer/_004_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens [3] ), .QN(\u2_ps2_cer/_065_ ) );
DFFR_X1 \u2_ps2_cer/_133_ ( .D(\u2_ps2_cer/_000_ ), .RN(clrn ), .CK(clk ), .Q(\u2_ps2_cer/counted ), .QN(\u2_ps2_cer/_066_ ) );
NOR2_X4 \u3_seg_h_0/_43_ ( .A1(\u3_seg_h_0/_31_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_01_ ) );
INV_X2 \u3_seg_h_0/_44_ ( .A(\u3_seg_h_0/_01_ ), .ZN(\u3_seg_h_0/_02_ ) );
INV_X4 \u3_seg_h_0/_45_ ( .A(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_03_ ) );
NOR2_X2 \u3_seg_h_0/_46_ ( .A1(\u3_seg_h_0/_03_ ), .A2(\u3_seg_h_0/_34_ ), .ZN(\u3_seg_h_0/_04_ ) );
INV_X16 \u3_seg_h_0/_47_ ( .A(\u3_seg_h_0/_34_ ), .ZN(\u3_seg_h_0/_05_ ) );
NOR2_X2 \u3_seg_h_0/_48_ ( .A1(\u3_seg_h_0/_05_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_06_ ) );
OR3_X4 \u3_seg_h_0/_49_ ( .A1(\u3_seg_h_0/_02_ ), .A2(\u3_seg_h_0/_04_ ), .A3(\u3_seg_h_0/_06_ ), .ZN(\u3_seg_h_0/_07_ ) );
INV_X32 \u3_seg_h_0/_50_ ( .A(\u3_seg_h_0/_31_ ), .ZN(\u3_seg_h_0/_08_ ) );
NOR2_X2 \u3_seg_h_0/_51_ ( .A1(\u3_seg_h_0/_08_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_09_ ) );
NOR2_X4 \u3_seg_h_0/_52_ ( .A1(\u3_seg_h_0/_34_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_10_ ) );
AND2_X1 \u3_seg_h_0/_53_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_10_ ), .ZN(\u3_seg_h_0/_11_ ) );
INV_X1 \u3_seg_h_0/_54_ ( .A(\u3_seg_h_0/_11_ ), .ZN(\u3_seg_h_0/_12_ ) );
INV_X1 \u3_seg_h_0/_55_ ( .A(\u3_seg_h_0/_00_ ), .ZN(\u3_seg_h_0/_13_ ) );
AND2_X4 \u3_seg_h_0/_56_ ( .A1(\u3_seg_h_0/_31_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_14_ ) );
AOI21_X1 \u3_seg_h_0/_57_ ( .A(\u3_seg_h_0/_13_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_15_ ) );
NAND3_X1 \u3_seg_h_0/_58_ ( .A1(\u3_seg_h_0/_07_ ), .A2(\u3_seg_h_0/_12_ ), .A3(\u3_seg_h_0/_15_ ), .ZN(\u3_seg_h_0/_35_ ) );
NAND2_X1 \u3_seg_h_0/_59_ ( .A1(\u3_seg_h_0/_02_ ), .A2(\u3_seg_h_0/_10_ ), .ZN(\u3_seg_h_0/_16_ ) );
AND2_X2 \u3_seg_h_0/_60_ ( .A1(\u3_seg_h_0/_34_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_17_ ) );
NAND2_X1 \u3_seg_h_0/_61_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_17_ ), .ZN(\u3_seg_h_0/_18_ ) );
NAND3_X1 \u3_seg_h_0/_62_ ( .A1(\u3_seg_h_0/_15_ ), .A2(\u3_seg_h_0/_16_ ), .A3(\u3_seg_h_0/_18_ ), .ZN(\u3_seg_h_0/_36_ ) );
NOR3_X1 \u3_seg_h_0/_63_ ( .A1(\u3_seg_h_0/_03_ ), .A2(\u3_seg_h_0/_34_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_19_ ) );
AOI21_X1 \u3_seg_h_0/_64_ ( .A(\u3_seg_h_0/_19_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_20_ ) );
NAND3_X1 \u3_seg_h_0/_65_ ( .A1(\u3_seg_h_0/_05_ ), .A2(\u3_seg_h_0/_03_ ), .A3(\u3_seg_h_0/_31_ ), .ZN(\u3_seg_h_0/_21_ ) );
NAND2_X1 \u3_seg_h_0/_66_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_06_ ), .ZN(\u3_seg_h_0/_22_ ) );
NAND4_X1 \u3_seg_h_0/_67_ ( .A1(\u3_seg_h_0/_20_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_21_ ), .A4(\u3_seg_h_0/_22_ ), .ZN(\u3_seg_h_0/_37_ ) );
NAND3_X1 \u3_seg_h_0/_68_ ( .A1(\u3_seg_h_0/_06_ ), .A2(\u3_seg_h_0/_08_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_23_ ) );
AOI22_X1 \u3_seg_h_0/_69_ ( .A1(\u3_seg_h_0/_04_ ), .A2(\u3_seg_h_0/_01_ ), .B1(\u3_seg_h_0/_14_ ), .B2(\u3_seg_h_0/_17_ ), .ZN(\u3_seg_h_0/_24_ ) );
NAND4_X1 \u3_seg_h_0/_70_ ( .A1(\u3_seg_h_0/_12_ ), .A2(\u3_seg_h_0/_15_ ), .A3(\u3_seg_h_0/_23_ ), .A4(\u3_seg_h_0/_24_ ), .ZN(\u3_seg_h_0/_38_ ) );
OAI21_X1 \u3_seg_h_0/_71_ ( .A(\u3_seg_h_0/_17_ ), .B1(\u3_seg_h_0/_08_ ), .B2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_25_ ) );
NAND3_X1 \u3_seg_h_0/_72_ ( .A1(\u3_seg_h_0/_10_ ), .A2(\u3_seg_h_0/_08_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_26_ ) );
NAND3_X1 \u3_seg_h_0/_73_ ( .A1(\u3_seg_h_0/_25_ ), .A2(\u3_seg_h_0/_26_ ), .A3(\u3_seg_h_0/_00_ ), .ZN(\u3_seg_h_0/_39_ ) );
AND2_X1 \u3_seg_h_0/_74_ ( .A1(\u3_seg_h_0/_08_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_27_ ) );
OAI21_X1 \u3_seg_h_0/_75_ ( .A(\u3_seg_h_0/_04_ ), .B1(\u3_seg_h_0/_27_ ), .B2(\u3_seg_h_0/_09_ ), .ZN(\u3_seg_h_0/_28_ ) );
NAND2_X1 \u3_seg_h_0/_76_ ( .A1(\u3_seg_h_0/_06_ ), .A2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_29_ ) );
NAND4_X1 \u3_seg_h_0/_77_ ( .A1(\u3_seg_h_0/_28_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_25_ ), .A4(\u3_seg_h_0/_29_ ), .ZN(\u3_seg_h_0/_40_ ) );
AOI22_X1 \u3_seg_h_0/_78_ ( .A1(\u3_seg_h_0/_10_ ), .A2(\u3_seg_h_0/_09_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_01_ ), .ZN(\u3_seg_h_0/_30_ ) );
NAND4_X1 \u3_seg_h_0/_79_ ( .A1(\u3_seg_h_0/_30_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_18_ ), .A4(\u3_seg_h_0/_29_ ), .ZN(\u3_seg_h_0/_41_ ) );
LOGIC1_X1 \u3_seg_h_0/_80_ ( .Z(\u3_seg_h_0/_42_ ) );
BUF_X1 \u3_seg_h_0/_81_ ( .A(\u3_seg_h_0/_42_ ), .Z(\seg_out_2 [0] ) );
BUF_X1 \u3_seg_h_0/_82_ ( .A(\key_ascii_display [3] ), .Z(\u3_seg_h_0/_34_ ) );
BUF_X1 \u3_seg_h_0/_83_ ( .A(\key_ascii_display [2] ), .Z(\u3_seg_h_0/_33_ ) );
BUF_X1 \u3_seg_h_0/_84_ ( .A(\key_ascii_display [0] ), .Z(\u3_seg_h_0/_31_ ) );
BUF_X1 \u3_seg_h_0/_85_ ( .A(\key_ascii_display [1] ), .Z(\u3_seg_h_0/_32_ ) );
BUF_X1 \u3_seg_h_0/_86_ ( .A(en ), .Z(\u3_seg_h_0/_00_ ) );
BUF_X1 \u3_seg_h_0/_87_ ( .A(\u3_seg_h_0/_35_ ), .Z(\seg_out_2 [1] ) );
BUF_X1 \u3_seg_h_0/_88_ ( .A(\u3_seg_h_0/_36_ ), .Z(\seg_out_2 [2] ) );
BUF_X1 \u3_seg_h_0/_89_ ( .A(\u3_seg_h_0/_37_ ), .Z(\seg_out_2 [3] ) );
BUF_X1 \u3_seg_h_0/_90_ ( .A(\u3_seg_h_0/_38_ ), .Z(\seg_out_2 [4] ) );
BUF_X1 \u3_seg_h_0/_91_ ( .A(\u3_seg_h_0/_39_ ), .Z(\seg_out_2 [5] ) );
BUF_X1 \u3_seg_h_0/_92_ ( .A(\u3_seg_h_0/_40_ ), .Z(\seg_out_2 [6] ) );
BUF_X1 \u3_seg_h_0/_93_ ( .A(\u3_seg_h_0/_41_ ), .Z(\seg_out_2 [7] ) );
NOR2_X4 \u4_seg_h_1/_43_ ( .A1(\u4_seg_h_1/_31_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_01_ ) );
INV_X2 \u4_seg_h_1/_44_ ( .A(\u4_seg_h_1/_01_ ), .ZN(\u4_seg_h_1/_02_ ) );
INV_X4 \u4_seg_h_1/_45_ ( .A(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_03_ ) );
NOR2_X2 \u4_seg_h_1/_46_ ( .A1(\u4_seg_h_1/_03_ ), .A2(\u4_seg_h_1/_34_ ), .ZN(\u4_seg_h_1/_04_ ) );
INV_X16 \u4_seg_h_1/_47_ ( .A(\u4_seg_h_1/_34_ ), .ZN(\u4_seg_h_1/_05_ ) );
NOR2_X2 \u4_seg_h_1/_48_ ( .A1(\u4_seg_h_1/_05_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_06_ ) );
OR3_X4 \u4_seg_h_1/_49_ ( .A1(\u4_seg_h_1/_02_ ), .A2(\u4_seg_h_1/_04_ ), .A3(\u4_seg_h_1/_06_ ), .ZN(\u4_seg_h_1/_07_ ) );
INV_X32 \u4_seg_h_1/_50_ ( .A(\u4_seg_h_1/_31_ ), .ZN(\u4_seg_h_1/_08_ ) );
NOR2_X2 \u4_seg_h_1/_51_ ( .A1(\u4_seg_h_1/_08_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_09_ ) );
NOR2_X4 \u4_seg_h_1/_52_ ( .A1(\u4_seg_h_1/_34_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_10_ ) );
AND2_X1 \u4_seg_h_1/_53_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_10_ ), .ZN(\u4_seg_h_1/_11_ ) );
INV_X1 \u4_seg_h_1/_54_ ( .A(\u4_seg_h_1/_11_ ), .ZN(\u4_seg_h_1/_12_ ) );
INV_X1 \u4_seg_h_1/_55_ ( .A(\u4_seg_h_1/_00_ ), .ZN(\u4_seg_h_1/_13_ ) );
AND2_X4 \u4_seg_h_1/_56_ ( .A1(\u4_seg_h_1/_31_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_14_ ) );
AOI21_X1 \u4_seg_h_1/_57_ ( .A(\u4_seg_h_1/_13_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_15_ ) );
NAND3_X1 \u4_seg_h_1/_58_ ( .A1(\u4_seg_h_1/_07_ ), .A2(\u4_seg_h_1/_12_ ), .A3(\u4_seg_h_1/_15_ ), .ZN(\u4_seg_h_1/_35_ ) );
NAND2_X1 \u4_seg_h_1/_59_ ( .A1(\u4_seg_h_1/_02_ ), .A2(\u4_seg_h_1/_10_ ), .ZN(\u4_seg_h_1/_16_ ) );
AND2_X2 \u4_seg_h_1/_60_ ( .A1(\u4_seg_h_1/_34_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_17_ ) );
NAND2_X1 \u4_seg_h_1/_61_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_17_ ), .ZN(\u4_seg_h_1/_18_ ) );
NAND3_X1 \u4_seg_h_1/_62_ ( .A1(\u4_seg_h_1/_15_ ), .A2(\u4_seg_h_1/_16_ ), .A3(\u4_seg_h_1/_18_ ), .ZN(\u4_seg_h_1/_36_ ) );
NOR3_X1 \u4_seg_h_1/_63_ ( .A1(\u4_seg_h_1/_03_ ), .A2(\u4_seg_h_1/_34_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_19_ ) );
AOI21_X1 \u4_seg_h_1/_64_ ( .A(\u4_seg_h_1/_19_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_20_ ) );
NAND3_X1 \u4_seg_h_1/_65_ ( .A1(\u4_seg_h_1/_05_ ), .A2(\u4_seg_h_1/_03_ ), .A3(\u4_seg_h_1/_31_ ), .ZN(\u4_seg_h_1/_21_ ) );
NAND2_X1 \u4_seg_h_1/_66_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_06_ ), .ZN(\u4_seg_h_1/_22_ ) );
NAND4_X1 \u4_seg_h_1/_67_ ( .A1(\u4_seg_h_1/_20_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_21_ ), .A4(\u4_seg_h_1/_22_ ), .ZN(\u4_seg_h_1/_37_ ) );
NAND3_X1 \u4_seg_h_1/_68_ ( .A1(\u4_seg_h_1/_06_ ), .A2(\u4_seg_h_1/_08_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_23_ ) );
AOI22_X1 \u4_seg_h_1/_69_ ( .A1(\u4_seg_h_1/_04_ ), .A2(\u4_seg_h_1/_01_ ), .B1(\u4_seg_h_1/_14_ ), .B2(\u4_seg_h_1/_17_ ), .ZN(\u4_seg_h_1/_24_ ) );
NAND4_X1 \u4_seg_h_1/_70_ ( .A1(\u4_seg_h_1/_12_ ), .A2(\u4_seg_h_1/_15_ ), .A3(\u4_seg_h_1/_23_ ), .A4(\u4_seg_h_1/_24_ ), .ZN(\u4_seg_h_1/_38_ ) );
OAI21_X1 \u4_seg_h_1/_71_ ( .A(\u4_seg_h_1/_17_ ), .B1(\u4_seg_h_1/_08_ ), .B2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_25_ ) );
NAND3_X1 \u4_seg_h_1/_72_ ( .A1(\u4_seg_h_1/_10_ ), .A2(\u4_seg_h_1/_08_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_26_ ) );
NAND3_X1 \u4_seg_h_1/_73_ ( .A1(\u4_seg_h_1/_25_ ), .A2(\u4_seg_h_1/_26_ ), .A3(\u4_seg_h_1/_00_ ), .ZN(\u4_seg_h_1/_39_ ) );
AND2_X1 \u4_seg_h_1/_74_ ( .A1(\u4_seg_h_1/_08_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_27_ ) );
OAI21_X1 \u4_seg_h_1/_75_ ( .A(\u4_seg_h_1/_04_ ), .B1(\u4_seg_h_1/_27_ ), .B2(\u4_seg_h_1/_09_ ), .ZN(\u4_seg_h_1/_28_ ) );
NAND2_X1 \u4_seg_h_1/_76_ ( .A1(\u4_seg_h_1/_06_ ), .A2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_29_ ) );
NAND4_X1 \u4_seg_h_1/_77_ ( .A1(\u4_seg_h_1/_28_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_25_ ), .A4(\u4_seg_h_1/_29_ ), .ZN(\u4_seg_h_1/_40_ ) );
AOI22_X1 \u4_seg_h_1/_78_ ( .A1(\u4_seg_h_1/_10_ ), .A2(\u4_seg_h_1/_09_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_01_ ), .ZN(\u4_seg_h_1/_30_ ) );
NAND4_X1 \u4_seg_h_1/_79_ ( .A1(\u4_seg_h_1/_30_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_18_ ), .A4(\u4_seg_h_1/_29_ ), .ZN(\u4_seg_h_1/_41_ ) );
LOGIC1_X1 \u4_seg_h_1/_80_ ( .Z(\u4_seg_h_1/_42_ ) );
BUF_X1 \u4_seg_h_1/_81_ ( .A(\u4_seg_h_1/_42_ ), .Z(\seg_out_3 [0] ) );
BUF_X1 \u4_seg_h_1/_82_ ( .A(\key_ascii_display [7] ), .Z(\u4_seg_h_1/_34_ ) );
BUF_X1 \u4_seg_h_1/_83_ ( .A(\key_ascii_display [6] ), .Z(\u4_seg_h_1/_33_ ) );
BUF_X1 \u4_seg_h_1/_84_ ( .A(\key_ascii_display [4] ), .Z(\u4_seg_h_1/_31_ ) );
BUF_X1 \u4_seg_h_1/_85_ ( .A(\key_ascii_display [5] ), .Z(\u4_seg_h_1/_32_ ) );
BUF_X1 \u4_seg_h_1/_86_ ( .A(en ), .Z(\u4_seg_h_1/_00_ ) );
BUF_X1 \u4_seg_h_1/_87_ ( .A(\u4_seg_h_1/_35_ ), .Z(\seg_out_3 [1] ) );
BUF_X1 \u4_seg_h_1/_88_ ( .A(\u4_seg_h_1/_36_ ), .Z(\seg_out_3 [2] ) );
BUF_X1 \u4_seg_h_1/_89_ ( .A(\u4_seg_h_1/_37_ ), .Z(\seg_out_3 [3] ) );
BUF_X1 \u4_seg_h_1/_90_ ( .A(\u4_seg_h_1/_38_ ), .Z(\seg_out_3 [4] ) );
BUF_X1 \u4_seg_h_1/_91_ ( .A(\u4_seg_h_1/_39_ ), .Z(\seg_out_3 [5] ) );
BUF_X1 \u4_seg_h_1/_92_ ( .A(\u4_seg_h_1/_40_ ), .Z(\seg_out_3 [6] ) );
BUF_X1 \u4_seg_h_1/_93_ ( .A(\u4_seg_h_1/_41_ ), .Z(\seg_out_3 [7] ) );
NOR2_X4 \u5_seg_h_2/_43_ ( .A1(\u5_seg_h_2/_31_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_01_ ) );
INV_X2 \u5_seg_h_2/_44_ ( .A(\u5_seg_h_2/_01_ ), .ZN(\u5_seg_h_2/_02_ ) );
INV_X4 \u5_seg_h_2/_45_ ( .A(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_03_ ) );
NOR2_X2 \u5_seg_h_2/_46_ ( .A1(\u5_seg_h_2/_03_ ), .A2(\u5_seg_h_2/_34_ ), .ZN(\u5_seg_h_2/_04_ ) );
INV_X16 \u5_seg_h_2/_47_ ( .A(\u5_seg_h_2/_34_ ), .ZN(\u5_seg_h_2/_05_ ) );
NOR2_X2 \u5_seg_h_2/_48_ ( .A1(\u5_seg_h_2/_05_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_06_ ) );
OR3_X4 \u5_seg_h_2/_49_ ( .A1(\u5_seg_h_2/_02_ ), .A2(\u5_seg_h_2/_04_ ), .A3(\u5_seg_h_2/_06_ ), .ZN(\u5_seg_h_2/_07_ ) );
INV_X32 \u5_seg_h_2/_50_ ( .A(\u5_seg_h_2/_31_ ), .ZN(\u5_seg_h_2/_08_ ) );
NOR2_X2 \u5_seg_h_2/_51_ ( .A1(\u5_seg_h_2/_08_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_09_ ) );
NOR2_X4 \u5_seg_h_2/_52_ ( .A1(\u5_seg_h_2/_34_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_10_ ) );
AND2_X1 \u5_seg_h_2/_53_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_10_ ), .ZN(\u5_seg_h_2/_11_ ) );
INV_X1 \u5_seg_h_2/_54_ ( .A(\u5_seg_h_2/_11_ ), .ZN(\u5_seg_h_2/_12_ ) );
INV_X1 \u5_seg_h_2/_55_ ( .A(\u5_seg_h_2/_00_ ), .ZN(\u5_seg_h_2/_13_ ) );
AND2_X4 \u5_seg_h_2/_56_ ( .A1(\u5_seg_h_2/_31_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_14_ ) );
AOI21_X1 \u5_seg_h_2/_57_ ( .A(\u5_seg_h_2/_13_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_15_ ) );
NAND3_X1 \u5_seg_h_2/_58_ ( .A1(\u5_seg_h_2/_07_ ), .A2(\u5_seg_h_2/_12_ ), .A3(\u5_seg_h_2/_15_ ), .ZN(\u5_seg_h_2/_35_ ) );
NAND2_X1 \u5_seg_h_2/_59_ ( .A1(\u5_seg_h_2/_02_ ), .A2(\u5_seg_h_2/_10_ ), .ZN(\u5_seg_h_2/_16_ ) );
AND2_X2 \u5_seg_h_2/_60_ ( .A1(\u5_seg_h_2/_34_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_17_ ) );
NAND2_X1 \u5_seg_h_2/_61_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_17_ ), .ZN(\u5_seg_h_2/_18_ ) );
NAND3_X1 \u5_seg_h_2/_62_ ( .A1(\u5_seg_h_2/_15_ ), .A2(\u5_seg_h_2/_16_ ), .A3(\u5_seg_h_2/_18_ ), .ZN(\u5_seg_h_2/_36_ ) );
NOR3_X1 \u5_seg_h_2/_63_ ( .A1(\u5_seg_h_2/_03_ ), .A2(\u5_seg_h_2/_34_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_19_ ) );
AOI21_X1 \u5_seg_h_2/_64_ ( .A(\u5_seg_h_2/_19_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_20_ ) );
NAND3_X1 \u5_seg_h_2/_65_ ( .A1(\u5_seg_h_2/_05_ ), .A2(\u5_seg_h_2/_03_ ), .A3(\u5_seg_h_2/_31_ ), .ZN(\u5_seg_h_2/_21_ ) );
NAND2_X1 \u5_seg_h_2/_66_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_06_ ), .ZN(\u5_seg_h_2/_22_ ) );
NAND4_X1 \u5_seg_h_2/_67_ ( .A1(\u5_seg_h_2/_20_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_21_ ), .A4(\u5_seg_h_2/_22_ ), .ZN(\u5_seg_h_2/_37_ ) );
NAND3_X1 \u5_seg_h_2/_68_ ( .A1(\u5_seg_h_2/_06_ ), .A2(\u5_seg_h_2/_08_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_23_ ) );
AOI22_X1 \u5_seg_h_2/_69_ ( .A1(\u5_seg_h_2/_04_ ), .A2(\u5_seg_h_2/_01_ ), .B1(\u5_seg_h_2/_14_ ), .B2(\u5_seg_h_2/_17_ ), .ZN(\u5_seg_h_2/_24_ ) );
NAND4_X1 \u5_seg_h_2/_70_ ( .A1(\u5_seg_h_2/_12_ ), .A2(\u5_seg_h_2/_15_ ), .A3(\u5_seg_h_2/_23_ ), .A4(\u5_seg_h_2/_24_ ), .ZN(\u5_seg_h_2/_38_ ) );
OAI21_X1 \u5_seg_h_2/_71_ ( .A(\u5_seg_h_2/_17_ ), .B1(\u5_seg_h_2/_08_ ), .B2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_25_ ) );
NAND3_X1 \u5_seg_h_2/_72_ ( .A1(\u5_seg_h_2/_10_ ), .A2(\u5_seg_h_2/_08_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_26_ ) );
NAND3_X1 \u5_seg_h_2/_73_ ( .A1(\u5_seg_h_2/_25_ ), .A2(\u5_seg_h_2/_26_ ), .A3(\u5_seg_h_2/_00_ ), .ZN(\u5_seg_h_2/_39_ ) );
AND2_X1 \u5_seg_h_2/_74_ ( .A1(\u5_seg_h_2/_08_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_27_ ) );
OAI21_X1 \u5_seg_h_2/_75_ ( .A(\u5_seg_h_2/_04_ ), .B1(\u5_seg_h_2/_27_ ), .B2(\u5_seg_h_2/_09_ ), .ZN(\u5_seg_h_2/_28_ ) );
NAND2_X1 \u5_seg_h_2/_76_ ( .A1(\u5_seg_h_2/_06_ ), .A2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_29_ ) );
NAND4_X1 \u5_seg_h_2/_77_ ( .A1(\u5_seg_h_2/_28_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_25_ ), .A4(\u5_seg_h_2/_29_ ), .ZN(\u5_seg_h_2/_40_ ) );
AOI22_X1 \u5_seg_h_2/_78_ ( .A1(\u5_seg_h_2/_10_ ), .A2(\u5_seg_h_2/_09_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_01_ ), .ZN(\u5_seg_h_2/_30_ ) );
NAND4_X1 \u5_seg_h_2/_79_ ( .A1(\u5_seg_h_2/_30_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_18_ ), .A4(\u5_seg_h_2/_29_ ), .ZN(\u5_seg_h_2/_41_ ) );
LOGIC1_X1 \u5_seg_h_2/_80_ ( .Z(\u5_seg_h_2/_42_ ) );
BUF_X1 \u5_seg_h_2/_81_ ( .A(\u5_seg_h_2/_42_ ), .Z(\seg_out_0 [0] ) );
BUF_X1 \u5_seg_h_2/_82_ ( .A(\key_scan_display [3] ), .Z(\u5_seg_h_2/_34_ ) );
BUF_X1 \u5_seg_h_2/_83_ ( .A(\key_scan_display [2] ), .Z(\u5_seg_h_2/_33_ ) );
BUF_X1 \u5_seg_h_2/_84_ ( .A(\key_scan_display [0] ), .Z(\u5_seg_h_2/_31_ ) );
BUF_X1 \u5_seg_h_2/_85_ ( .A(\key_scan_display [1] ), .Z(\u5_seg_h_2/_32_ ) );
BUF_X1 \u5_seg_h_2/_86_ ( .A(en ), .Z(\u5_seg_h_2/_00_ ) );
BUF_X1 \u5_seg_h_2/_87_ ( .A(\u5_seg_h_2/_35_ ), .Z(\seg_out_0 [1] ) );
BUF_X1 \u5_seg_h_2/_88_ ( .A(\u5_seg_h_2/_36_ ), .Z(\seg_out_0 [2] ) );
BUF_X1 \u5_seg_h_2/_89_ ( .A(\u5_seg_h_2/_37_ ), .Z(\seg_out_0 [3] ) );
BUF_X1 \u5_seg_h_2/_90_ ( .A(\u5_seg_h_2/_38_ ), .Z(\seg_out_0 [4] ) );
BUF_X1 \u5_seg_h_2/_91_ ( .A(\u5_seg_h_2/_39_ ), .Z(\seg_out_0 [5] ) );
BUF_X1 \u5_seg_h_2/_92_ ( .A(\u5_seg_h_2/_40_ ), .Z(\seg_out_0 [6] ) );
BUF_X1 \u5_seg_h_2/_93_ ( .A(\u5_seg_h_2/_41_ ), .Z(\seg_out_0 [7] ) );
NOR2_X4 \u6_seg_h_3/_43_ ( .A1(\u6_seg_h_3/_31_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_01_ ) );
INV_X2 \u6_seg_h_3/_44_ ( .A(\u6_seg_h_3/_01_ ), .ZN(\u6_seg_h_3/_02_ ) );
INV_X4 \u6_seg_h_3/_45_ ( .A(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_03_ ) );
NOR2_X2 \u6_seg_h_3/_46_ ( .A1(\u6_seg_h_3/_03_ ), .A2(\u6_seg_h_3/_34_ ), .ZN(\u6_seg_h_3/_04_ ) );
INV_X16 \u6_seg_h_3/_47_ ( .A(\u6_seg_h_3/_34_ ), .ZN(\u6_seg_h_3/_05_ ) );
NOR2_X2 \u6_seg_h_3/_48_ ( .A1(\u6_seg_h_3/_05_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_06_ ) );
OR3_X4 \u6_seg_h_3/_49_ ( .A1(\u6_seg_h_3/_02_ ), .A2(\u6_seg_h_3/_04_ ), .A3(\u6_seg_h_3/_06_ ), .ZN(\u6_seg_h_3/_07_ ) );
INV_X32 \u6_seg_h_3/_50_ ( .A(\u6_seg_h_3/_31_ ), .ZN(\u6_seg_h_3/_08_ ) );
NOR2_X2 \u6_seg_h_3/_51_ ( .A1(\u6_seg_h_3/_08_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_09_ ) );
NOR2_X4 \u6_seg_h_3/_52_ ( .A1(\u6_seg_h_3/_34_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_10_ ) );
AND2_X1 \u6_seg_h_3/_53_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_10_ ), .ZN(\u6_seg_h_3/_11_ ) );
INV_X1 \u6_seg_h_3/_54_ ( .A(\u6_seg_h_3/_11_ ), .ZN(\u6_seg_h_3/_12_ ) );
INV_X1 \u6_seg_h_3/_55_ ( .A(\u6_seg_h_3/_00_ ), .ZN(\u6_seg_h_3/_13_ ) );
AND2_X4 \u6_seg_h_3/_56_ ( .A1(\u6_seg_h_3/_31_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_14_ ) );
AOI21_X1 \u6_seg_h_3/_57_ ( .A(\u6_seg_h_3/_13_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_15_ ) );
NAND3_X1 \u6_seg_h_3/_58_ ( .A1(\u6_seg_h_3/_07_ ), .A2(\u6_seg_h_3/_12_ ), .A3(\u6_seg_h_3/_15_ ), .ZN(\u6_seg_h_3/_35_ ) );
NAND2_X1 \u6_seg_h_3/_59_ ( .A1(\u6_seg_h_3/_02_ ), .A2(\u6_seg_h_3/_10_ ), .ZN(\u6_seg_h_3/_16_ ) );
AND2_X2 \u6_seg_h_3/_60_ ( .A1(\u6_seg_h_3/_34_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_17_ ) );
NAND2_X1 \u6_seg_h_3/_61_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_17_ ), .ZN(\u6_seg_h_3/_18_ ) );
NAND3_X1 \u6_seg_h_3/_62_ ( .A1(\u6_seg_h_3/_15_ ), .A2(\u6_seg_h_3/_16_ ), .A3(\u6_seg_h_3/_18_ ), .ZN(\u6_seg_h_3/_36_ ) );
NOR3_X1 \u6_seg_h_3/_63_ ( .A1(\u6_seg_h_3/_03_ ), .A2(\u6_seg_h_3/_34_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_19_ ) );
AOI21_X1 \u6_seg_h_3/_64_ ( .A(\u6_seg_h_3/_19_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_20_ ) );
NAND3_X1 \u6_seg_h_3/_65_ ( .A1(\u6_seg_h_3/_05_ ), .A2(\u6_seg_h_3/_03_ ), .A3(\u6_seg_h_3/_31_ ), .ZN(\u6_seg_h_3/_21_ ) );
NAND2_X1 \u6_seg_h_3/_66_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_06_ ), .ZN(\u6_seg_h_3/_22_ ) );
NAND4_X1 \u6_seg_h_3/_67_ ( .A1(\u6_seg_h_3/_20_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_21_ ), .A4(\u6_seg_h_3/_22_ ), .ZN(\u6_seg_h_3/_37_ ) );
NAND3_X1 \u6_seg_h_3/_68_ ( .A1(\u6_seg_h_3/_06_ ), .A2(\u6_seg_h_3/_08_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_23_ ) );
AOI22_X1 \u6_seg_h_3/_69_ ( .A1(\u6_seg_h_3/_04_ ), .A2(\u6_seg_h_3/_01_ ), .B1(\u6_seg_h_3/_14_ ), .B2(\u6_seg_h_3/_17_ ), .ZN(\u6_seg_h_3/_24_ ) );
NAND4_X1 \u6_seg_h_3/_70_ ( .A1(\u6_seg_h_3/_12_ ), .A2(\u6_seg_h_3/_15_ ), .A3(\u6_seg_h_3/_23_ ), .A4(\u6_seg_h_3/_24_ ), .ZN(\u6_seg_h_3/_38_ ) );
OAI21_X1 \u6_seg_h_3/_71_ ( .A(\u6_seg_h_3/_17_ ), .B1(\u6_seg_h_3/_08_ ), .B2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_25_ ) );
NAND3_X1 \u6_seg_h_3/_72_ ( .A1(\u6_seg_h_3/_10_ ), .A2(\u6_seg_h_3/_08_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_26_ ) );
NAND3_X1 \u6_seg_h_3/_73_ ( .A1(\u6_seg_h_3/_25_ ), .A2(\u6_seg_h_3/_26_ ), .A3(\u6_seg_h_3/_00_ ), .ZN(\u6_seg_h_3/_39_ ) );
AND2_X1 \u6_seg_h_3/_74_ ( .A1(\u6_seg_h_3/_08_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_27_ ) );
OAI21_X1 \u6_seg_h_3/_75_ ( .A(\u6_seg_h_3/_04_ ), .B1(\u6_seg_h_3/_27_ ), .B2(\u6_seg_h_3/_09_ ), .ZN(\u6_seg_h_3/_28_ ) );
NAND2_X1 \u6_seg_h_3/_76_ ( .A1(\u6_seg_h_3/_06_ ), .A2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_29_ ) );
NAND4_X1 \u6_seg_h_3/_77_ ( .A1(\u6_seg_h_3/_28_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_25_ ), .A4(\u6_seg_h_3/_29_ ), .ZN(\u6_seg_h_3/_40_ ) );
AOI22_X1 \u6_seg_h_3/_78_ ( .A1(\u6_seg_h_3/_10_ ), .A2(\u6_seg_h_3/_09_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_01_ ), .ZN(\u6_seg_h_3/_30_ ) );
NAND4_X1 \u6_seg_h_3/_79_ ( .A1(\u6_seg_h_3/_30_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_18_ ), .A4(\u6_seg_h_3/_29_ ), .ZN(\u6_seg_h_3/_41_ ) );
LOGIC1_X1 \u6_seg_h_3/_80_ ( .Z(\u6_seg_h_3/_42_ ) );
BUF_X1 \u6_seg_h_3/_81_ ( .A(\u6_seg_h_3/_42_ ), .Z(\seg_out_1 [0] ) );
BUF_X1 \u6_seg_h_3/_82_ ( .A(\key_scan_display [7] ), .Z(\u6_seg_h_3/_34_ ) );
BUF_X1 \u6_seg_h_3/_83_ ( .A(\key_scan_display [6] ), .Z(\u6_seg_h_3/_33_ ) );
BUF_X1 \u6_seg_h_3/_84_ ( .A(\key_scan_display [4] ), .Z(\u6_seg_h_3/_31_ ) );
BUF_X1 \u6_seg_h_3/_85_ ( .A(\key_scan_display [5] ), .Z(\u6_seg_h_3/_32_ ) );
BUF_X1 \u6_seg_h_3/_86_ ( .A(en ), .Z(\u6_seg_h_3/_00_ ) );
BUF_X1 \u6_seg_h_3/_87_ ( .A(\u6_seg_h_3/_35_ ), .Z(\seg_out_1 [1] ) );
BUF_X1 \u6_seg_h_3/_88_ ( .A(\u6_seg_h_3/_36_ ), .Z(\seg_out_1 [2] ) );
BUF_X1 \u6_seg_h_3/_89_ ( .A(\u6_seg_h_3/_37_ ), .Z(\seg_out_1 [3] ) );
BUF_X1 \u6_seg_h_3/_90_ ( .A(\u6_seg_h_3/_38_ ), .Z(\seg_out_1 [4] ) );
BUF_X1 \u6_seg_h_3/_91_ ( .A(\u6_seg_h_3/_39_ ), .Z(\seg_out_1 [5] ) );
BUF_X1 \u6_seg_h_3/_92_ ( .A(\u6_seg_h_3/_40_ ), .Z(\seg_out_1 [6] ) );
BUF_X1 \u6_seg_h_3/_93_ ( .A(\u6_seg_h_3/_41_ ), .Z(\seg_out_1 [7] ) );
NOR2_X4 \u7_seg_h_4/_43_ ( .A1(\u7_seg_h_4/_31_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_01_ ) );
INV_X2 \u7_seg_h_4/_44_ ( .A(\u7_seg_h_4/_01_ ), .ZN(\u7_seg_h_4/_02_ ) );
INV_X4 \u7_seg_h_4/_45_ ( .A(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_03_ ) );
NOR2_X2 \u7_seg_h_4/_46_ ( .A1(\u7_seg_h_4/_03_ ), .A2(\u7_seg_h_4/_34_ ), .ZN(\u7_seg_h_4/_04_ ) );
INV_X16 \u7_seg_h_4/_47_ ( .A(\u7_seg_h_4/_34_ ), .ZN(\u7_seg_h_4/_05_ ) );
NOR2_X2 \u7_seg_h_4/_48_ ( .A1(\u7_seg_h_4/_05_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_06_ ) );
OR3_X4 \u7_seg_h_4/_49_ ( .A1(\u7_seg_h_4/_02_ ), .A2(\u7_seg_h_4/_04_ ), .A3(\u7_seg_h_4/_06_ ), .ZN(\u7_seg_h_4/_07_ ) );
INV_X32 \u7_seg_h_4/_50_ ( .A(\u7_seg_h_4/_31_ ), .ZN(\u7_seg_h_4/_08_ ) );
NOR2_X2 \u7_seg_h_4/_51_ ( .A1(\u7_seg_h_4/_08_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_09_ ) );
NOR2_X4 \u7_seg_h_4/_52_ ( .A1(\u7_seg_h_4/_34_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_10_ ) );
AND2_X1 \u7_seg_h_4/_53_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_10_ ), .ZN(\u7_seg_h_4/_11_ ) );
INV_X1 \u7_seg_h_4/_54_ ( .A(\u7_seg_h_4/_11_ ), .ZN(\u7_seg_h_4/_12_ ) );
INV_X1 \u7_seg_h_4/_55_ ( .A(\u7_seg_h_4/_00_ ), .ZN(\u7_seg_h_4/_13_ ) );
AND2_X4 \u7_seg_h_4/_56_ ( .A1(\u7_seg_h_4/_31_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_14_ ) );
AOI21_X1 \u7_seg_h_4/_57_ ( .A(\u7_seg_h_4/_13_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_15_ ) );
NAND3_X1 \u7_seg_h_4/_58_ ( .A1(\u7_seg_h_4/_07_ ), .A2(\u7_seg_h_4/_12_ ), .A3(\u7_seg_h_4/_15_ ), .ZN(\u7_seg_h_4/_35_ ) );
NAND2_X1 \u7_seg_h_4/_59_ ( .A1(\u7_seg_h_4/_02_ ), .A2(\u7_seg_h_4/_10_ ), .ZN(\u7_seg_h_4/_16_ ) );
AND2_X2 \u7_seg_h_4/_60_ ( .A1(\u7_seg_h_4/_34_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_17_ ) );
NAND2_X1 \u7_seg_h_4/_61_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_17_ ), .ZN(\u7_seg_h_4/_18_ ) );
NAND3_X1 \u7_seg_h_4/_62_ ( .A1(\u7_seg_h_4/_15_ ), .A2(\u7_seg_h_4/_16_ ), .A3(\u7_seg_h_4/_18_ ), .ZN(\u7_seg_h_4/_36_ ) );
NOR3_X1 \u7_seg_h_4/_63_ ( .A1(\u7_seg_h_4/_03_ ), .A2(\u7_seg_h_4/_34_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_19_ ) );
AOI21_X1 \u7_seg_h_4/_64_ ( .A(\u7_seg_h_4/_19_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_20_ ) );
NAND3_X1 \u7_seg_h_4/_65_ ( .A1(\u7_seg_h_4/_05_ ), .A2(\u7_seg_h_4/_03_ ), .A3(\u7_seg_h_4/_31_ ), .ZN(\u7_seg_h_4/_21_ ) );
NAND2_X1 \u7_seg_h_4/_66_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_06_ ), .ZN(\u7_seg_h_4/_22_ ) );
NAND4_X1 \u7_seg_h_4/_67_ ( .A1(\u7_seg_h_4/_20_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_21_ ), .A4(\u7_seg_h_4/_22_ ), .ZN(\u7_seg_h_4/_37_ ) );
NAND3_X1 \u7_seg_h_4/_68_ ( .A1(\u7_seg_h_4/_06_ ), .A2(\u7_seg_h_4/_08_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_23_ ) );
AOI22_X1 \u7_seg_h_4/_69_ ( .A1(\u7_seg_h_4/_04_ ), .A2(\u7_seg_h_4/_01_ ), .B1(\u7_seg_h_4/_14_ ), .B2(\u7_seg_h_4/_17_ ), .ZN(\u7_seg_h_4/_24_ ) );
NAND4_X1 \u7_seg_h_4/_70_ ( .A1(\u7_seg_h_4/_12_ ), .A2(\u7_seg_h_4/_15_ ), .A3(\u7_seg_h_4/_23_ ), .A4(\u7_seg_h_4/_24_ ), .ZN(\u7_seg_h_4/_38_ ) );
OAI21_X1 \u7_seg_h_4/_71_ ( .A(\u7_seg_h_4/_17_ ), .B1(\u7_seg_h_4/_08_ ), .B2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_25_ ) );
NAND3_X1 \u7_seg_h_4/_72_ ( .A1(\u7_seg_h_4/_10_ ), .A2(\u7_seg_h_4/_08_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_26_ ) );
NAND3_X1 \u7_seg_h_4/_73_ ( .A1(\u7_seg_h_4/_25_ ), .A2(\u7_seg_h_4/_26_ ), .A3(\u7_seg_h_4/_00_ ), .ZN(\u7_seg_h_4/_39_ ) );
AND2_X1 \u7_seg_h_4/_74_ ( .A1(\u7_seg_h_4/_08_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_27_ ) );
OAI21_X1 \u7_seg_h_4/_75_ ( .A(\u7_seg_h_4/_04_ ), .B1(\u7_seg_h_4/_27_ ), .B2(\u7_seg_h_4/_09_ ), .ZN(\u7_seg_h_4/_28_ ) );
NAND2_X1 \u7_seg_h_4/_76_ ( .A1(\u7_seg_h_4/_06_ ), .A2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_29_ ) );
NAND4_X1 \u7_seg_h_4/_77_ ( .A1(\u7_seg_h_4/_28_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_25_ ), .A4(\u7_seg_h_4/_29_ ), .ZN(\u7_seg_h_4/_40_ ) );
AOI22_X1 \u7_seg_h_4/_78_ ( .A1(\u7_seg_h_4/_10_ ), .A2(\u7_seg_h_4/_09_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_01_ ), .ZN(\u7_seg_h_4/_30_ ) );
NAND4_X1 \u7_seg_h_4/_79_ ( .A1(\u7_seg_h_4/_30_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_18_ ), .A4(\u7_seg_h_4/_29_ ), .ZN(\u7_seg_h_4/_41_ ) );
LOGIC1_X1 \u7_seg_h_4/_80_ ( .Z(\u7_seg_h_4/_42_ ) );
BUF_X1 \u7_seg_h_4/_81_ ( .A(\u7_seg_h_4/_42_ ), .Z(\seg_out_4 [0] ) );
BUF_X1 \u7_seg_h_4/_82_ ( .A(\high_units [3] ), .Z(\u7_seg_h_4/_34_ ) );
BUF_X1 \u7_seg_h_4/_83_ ( .A(\high_units [2] ), .Z(\u7_seg_h_4/_33_ ) );
BUF_X1 \u7_seg_h_4/_84_ ( .A(\high_units [0] ), .Z(\u7_seg_h_4/_31_ ) );
BUF_X1 \u7_seg_h_4/_85_ ( .A(\high_units [1] ), .Z(\u7_seg_h_4/_32_ ) );
BUF_X1 \u7_seg_h_4/_86_ ( .A(_132_ ), .Z(\u7_seg_h_4/_00_ ) );
BUF_X1 \u7_seg_h_4/_87_ ( .A(\u7_seg_h_4/_35_ ), .Z(\seg_out_4 [1] ) );
BUF_X1 \u7_seg_h_4/_88_ ( .A(\u7_seg_h_4/_36_ ), .Z(\seg_out_4 [2] ) );
BUF_X1 \u7_seg_h_4/_89_ ( .A(\u7_seg_h_4/_37_ ), .Z(\seg_out_4 [3] ) );
BUF_X1 \u7_seg_h_4/_90_ ( .A(\u7_seg_h_4/_38_ ), .Z(\seg_out_4 [4] ) );
BUF_X1 \u7_seg_h_4/_91_ ( .A(\u7_seg_h_4/_39_ ), .Z(\seg_out_4 [5] ) );
BUF_X1 \u7_seg_h_4/_92_ ( .A(\u7_seg_h_4/_40_ ), .Z(\seg_out_4 [6] ) );
BUF_X1 \u7_seg_h_4/_93_ ( .A(\u7_seg_h_4/_41_ ), .Z(\seg_out_4 [7] ) );
NOR2_X4 \u8_seg_h_5/_43_ ( .A1(\u8_seg_h_5/_31_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_01_ ) );
INV_X2 \u8_seg_h_5/_44_ ( .A(\u8_seg_h_5/_01_ ), .ZN(\u8_seg_h_5/_02_ ) );
INV_X4 \u8_seg_h_5/_45_ ( .A(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_03_ ) );
NOR2_X2 \u8_seg_h_5/_46_ ( .A1(\u8_seg_h_5/_03_ ), .A2(\u8_seg_h_5/_34_ ), .ZN(\u8_seg_h_5/_04_ ) );
INV_X16 \u8_seg_h_5/_47_ ( .A(\u8_seg_h_5/_34_ ), .ZN(\u8_seg_h_5/_05_ ) );
NOR2_X2 \u8_seg_h_5/_48_ ( .A1(\u8_seg_h_5/_05_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_06_ ) );
OR3_X4 \u8_seg_h_5/_49_ ( .A1(\u8_seg_h_5/_02_ ), .A2(\u8_seg_h_5/_04_ ), .A3(\u8_seg_h_5/_06_ ), .ZN(\u8_seg_h_5/_07_ ) );
INV_X32 \u8_seg_h_5/_50_ ( .A(\u8_seg_h_5/_31_ ), .ZN(\u8_seg_h_5/_08_ ) );
NOR2_X2 \u8_seg_h_5/_51_ ( .A1(\u8_seg_h_5/_08_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_09_ ) );
NOR2_X4 \u8_seg_h_5/_52_ ( .A1(\u8_seg_h_5/_34_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_10_ ) );
AND2_X1 \u8_seg_h_5/_53_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_10_ ), .ZN(\u8_seg_h_5/_11_ ) );
INV_X1 \u8_seg_h_5/_54_ ( .A(\u8_seg_h_5/_11_ ), .ZN(\u8_seg_h_5/_12_ ) );
INV_X1 \u8_seg_h_5/_55_ ( .A(\u8_seg_h_5/_00_ ), .ZN(\u8_seg_h_5/_13_ ) );
AND2_X4 \u8_seg_h_5/_56_ ( .A1(\u8_seg_h_5/_31_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_14_ ) );
AOI21_X1 \u8_seg_h_5/_57_ ( .A(\u8_seg_h_5/_13_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_15_ ) );
NAND3_X1 \u8_seg_h_5/_58_ ( .A1(\u8_seg_h_5/_07_ ), .A2(\u8_seg_h_5/_12_ ), .A3(\u8_seg_h_5/_15_ ), .ZN(\u8_seg_h_5/_35_ ) );
NAND2_X1 \u8_seg_h_5/_59_ ( .A1(\u8_seg_h_5/_02_ ), .A2(\u8_seg_h_5/_10_ ), .ZN(\u8_seg_h_5/_16_ ) );
AND2_X2 \u8_seg_h_5/_60_ ( .A1(\u8_seg_h_5/_34_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_17_ ) );
NAND2_X1 \u8_seg_h_5/_61_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_17_ ), .ZN(\u8_seg_h_5/_18_ ) );
NAND3_X1 \u8_seg_h_5/_62_ ( .A1(\u8_seg_h_5/_15_ ), .A2(\u8_seg_h_5/_16_ ), .A3(\u8_seg_h_5/_18_ ), .ZN(\u8_seg_h_5/_36_ ) );
NOR3_X1 \u8_seg_h_5/_63_ ( .A1(\u8_seg_h_5/_03_ ), .A2(\u8_seg_h_5/_34_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_19_ ) );
AOI21_X1 \u8_seg_h_5/_64_ ( .A(\u8_seg_h_5/_19_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_20_ ) );
NAND3_X1 \u8_seg_h_5/_65_ ( .A1(\u8_seg_h_5/_05_ ), .A2(\u8_seg_h_5/_03_ ), .A3(\u8_seg_h_5/_31_ ), .ZN(\u8_seg_h_5/_21_ ) );
NAND2_X1 \u8_seg_h_5/_66_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_06_ ), .ZN(\u8_seg_h_5/_22_ ) );
NAND4_X1 \u8_seg_h_5/_67_ ( .A1(\u8_seg_h_5/_20_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_21_ ), .A4(\u8_seg_h_5/_22_ ), .ZN(\u8_seg_h_5/_37_ ) );
NAND3_X1 \u8_seg_h_5/_68_ ( .A1(\u8_seg_h_5/_06_ ), .A2(\u8_seg_h_5/_08_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_23_ ) );
AOI22_X1 \u8_seg_h_5/_69_ ( .A1(\u8_seg_h_5/_04_ ), .A2(\u8_seg_h_5/_01_ ), .B1(\u8_seg_h_5/_14_ ), .B2(\u8_seg_h_5/_17_ ), .ZN(\u8_seg_h_5/_24_ ) );
NAND4_X1 \u8_seg_h_5/_70_ ( .A1(\u8_seg_h_5/_12_ ), .A2(\u8_seg_h_5/_15_ ), .A3(\u8_seg_h_5/_23_ ), .A4(\u8_seg_h_5/_24_ ), .ZN(\u8_seg_h_5/_38_ ) );
OAI21_X1 \u8_seg_h_5/_71_ ( .A(\u8_seg_h_5/_17_ ), .B1(\u8_seg_h_5/_08_ ), .B2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_25_ ) );
NAND3_X1 \u8_seg_h_5/_72_ ( .A1(\u8_seg_h_5/_10_ ), .A2(\u8_seg_h_5/_08_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_26_ ) );
NAND3_X1 \u8_seg_h_5/_73_ ( .A1(\u8_seg_h_5/_25_ ), .A2(\u8_seg_h_5/_26_ ), .A3(\u8_seg_h_5/_00_ ), .ZN(\u8_seg_h_5/_39_ ) );
AND2_X1 \u8_seg_h_5/_74_ ( .A1(\u8_seg_h_5/_08_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_27_ ) );
OAI21_X1 \u8_seg_h_5/_75_ ( .A(\u8_seg_h_5/_04_ ), .B1(\u8_seg_h_5/_27_ ), .B2(\u8_seg_h_5/_09_ ), .ZN(\u8_seg_h_5/_28_ ) );
NAND2_X1 \u8_seg_h_5/_76_ ( .A1(\u8_seg_h_5/_06_ ), .A2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_29_ ) );
NAND4_X1 \u8_seg_h_5/_77_ ( .A1(\u8_seg_h_5/_28_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_25_ ), .A4(\u8_seg_h_5/_29_ ), .ZN(\u8_seg_h_5/_40_ ) );
AOI22_X1 \u8_seg_h_5/_78_ ( .A1(\u8_seg_h_5/_10_ ), .A2(\u8_seg_h_5/_09_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_01_ ), .ZN(\u8_seg_h_5/_30_ ) );
NAND4_X1 \u8_seg_h_5/_79_ ( .A1(\u8_seg_h_5/_30_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_18_ ), .A4(\u8_seg_h_5/_29_ ), .ZN(\u8_seg_h_5/_41_ ) );
LOGIC1_X1 \u8_seg_h_5/_80_ ( .Z(\u8_seg_h_5/_42_ ) );
BUF_X1 \u8_seg_h_5/_81_ ( .A(\u8_seg_h_5/_42_ ), .Z(\seg_out_5 [0] ) );
BUF_X1 \u8_seg_h_5/_82_ ( .A(\high_tens [3] ), .Z(\u8_seg_h_5/_34_ ) );
BUF_X1 \u8_seg_h_5/_83_ ( .A(\high_tens [2] ), .Z(\u8_seg_h_5/_33_ ) );
BUF_X1 \u8_seg_h_5/_84_ ( .A(\high_tens [0] ), .Z(\u8_seg_h_5/_31_ ) );
BUF_X1 \u8_seg_h_5/_85_ ( .A(\high_tens [1] ), .Z(\u8_seg_h_5/_32_ ) );
BUF_X1 \u8_seg_h_5/_86_ ( .A(_132_ ), .Z(\u8_seg_h_5/_00_ ) );
BUF_X1 \u8_seg_h_5/_87_ ( .A(\u8_seg_h_5/_35_ ), .Z(\seg_out_5 [1] ) );
BUF_X1 \u8_seg_h_5/_88_ ( .A(\u8_seg_h_5/_36_ ), .Z(\seg_out_5 [2] ) );
BUF_X1 \u8_seg_h_5/_89_ ( .A(\u8_seg_h_5/_37_ ), .Z(\seg_out_5 [3] ) );
BUF_X1 \u8_seg_h_5/_90_ ( .A(\u8_seg_h_5/_38_ ), .Z(\seg_out_5 [4] ) );
BUF_X1 \u8_seg_h_5/_91_ ( .A(\u8_seg_h_5/_39_ ), .Z(\seg_out_5 [5] ) );
BUF_X1 \u8_seg_h_5/_92_ ( .A(\u8_seg_h_5/_40_ ), .Z(\seg_out_5 [6] ) );
BUF_X1 \u8_seg_h_5/_93_ ( .A(\u8_seg_h_5/_41_ ), .Z(\seg_out_5 [7] ) );
BUF_X8 fanout_buf_1 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\u1_ps2_dsh/_050_ ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\u1_ps2_dsh/_051_ ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\u1_ps2_dsh/key_ascii/i0/_0008_ ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\u1_ps2_dsh/key_ascii/i0/_0009_ ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\u1_ps2_dsh/key_ascii/i0/_0010_ ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\u1_ps2_dsh/key_ascii/i0/_0011_ ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\u1_ps2_dsh/key_ascii/i0/_0012_ ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\u1_ps2_dsh/key_ascii/i0/_0013_ ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\u1_ps2_dsh/key_ascii/i0/_0014_ ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\u1_ps2_dsh/key_ascii/i0/_0015_ ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(clrn ), .Z(fanout_net_28 ) );

endmodule
