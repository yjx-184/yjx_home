//Generate the verilog at 2024-12-03T15:15:21
module ps2_top (
clk,
clrn,
overflow,
ps2_clk,
ps2_data,
seg_out_0,
seg_out_1,
seg_out_2,
seg_out_3,
seg_out_4,
seg_out_5
);

input clk ;
input clrn ;
output overflow ;
input ps2_clk ;
input ps2_data ;
output [7:0] seg_out_0 ;
output [7:0] seg_out_1 ;
output [7:0] seg_out_2 ;
output [7:0] seg_out_3 ;
output [7:0] seg_out_4 ;
output [7:0] seg_out_5 ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire en ;
wire key_release ;
wire nextdata_n ;
wire ready ;
wire ready_d1 ;
wire \u0_ps2_kb/_0000_ ;
wire \u0_ps2_kb/_0001_ ;
wire \u0_ps2_kb/_0002_ ;
wire \u0_ps2_kb/_0003_ ;
wire \u0_ps2_kb/_0004_ ;
wire \u0_ps2_kb/_0005_ ;
wire \u0_ps2_kb/_0006_ ;
wire \u0_ps2_kb/_0007_ ;
wire \u0_ps2_kb/_0008_ ;
wire \u0_ps2_kb/_0009_ ;
wire \u0_ps2_kb/_0010_ ;
wire \u0_ps2_kb/_0011_ ;
wire \u0_ps2_kb/_0012_ ;
wire \u0_ps2_kb/_0013_ ;
wire \u0_ps2_kb/_0014_ ;
wire \u0_ps2_kb/_0015_ ;
wire \u0_ps2_kb/_0016_ ;
wire \u0_ps2_kb/_0017_ ;
wire \u0_ps2_kb/_0018_ ;
wire \u0_ps2_kb/_0019_ ;
wire \u0_ps2_kb/_0020_ ;
wire \u0_ps2_kb/_0021_ ;
wire \u0_ps2_kb/_0022_ ;
wire \u0_ps2_kb/_0023_ ;
wire \u0_ps2_kb/_0024_ ;
wire \u0_ps2_kb/_0025_ ;
wire \u0_ps2_kb/_0026_ ;
wire \u0_ps2_kb/_0027_ ;
wire \u0_ps2_kb/_0028_ ;
wire \u0_ps2_kb/_0029_ ;
wire \u0_ps2_kb/_0030_ ;
wire \u0_ps2_kb/_0031_ ;
wire \u0_ps2_kb/_0032_ ;
wire \u0_ps2_kb/_0033_ ;
wire \u0_ps2_kb/_0034_ ;
wire \u0_ps2_kb/_0035_ ;
wire \u0_ps2_kb/_0036_ ;
wire \u0_ps2_kb/_0037_ ;
wire \u0_ps2_kb/_0038_ ;
wire \u0_ps2_kb/_0039_ ;
wire \u0_ps2_kb/_0040_ ;
wire \u0_ps2_kb/_0041_ ;
wire \u0_ps2_kb/_0042_ ;
wire \u0_ps2_kb/_0043_ ;
wire \u0_ps2_kb/_0044_ ;
wire \u0_ps2_kb/_0045_ ;
wire \u0_ps2_kb/_0046_ ;
wire \u0_ps2_kb/_0047_ ;
wire \u0_ps2_kb/_0048_ ;
wire \u0_ps2_kb/_0049_ ;
wire \u0_ps2_kb/_0050_ ;
wire \u0_ps2_kb/_0051_ ;
wire \u0_ps2_kb/_0052_ ;
wire \u0_ps2_kb/_0053_ ;
wire \u0_ps2_kb/_0054_ ;
wire \u0_ps2_kb/_0055_ ;
wire \u0_ps2_kb/_0056_ ;
wire \u0_ps2_kb/_0057_ ;
wire \u0_ps2_kb/_0058_ ;
wire \u0_ps2_kb/_0059_ ;
wire \u0_ps2_kb/_0060_ ;
wire \u0_ps2_kb/_0061_ ;
wire \u0_ps2_kb/_0062_ ;
wire \u0_ps2_kb/_0063_ ;
wire \u0_ps2_kb/_0064_ ;
wire \u0_ps2_kb/_0065_ ;
wire \u0_ps2_kb/_0066_ ;
wire \u0_ps2_kb/_0067_ ;
wire \u0_ps2_kb/_0068_ ;
wire \u0_ps2_kb/_0069_ ;
wire \u0_ps2_kb/_0070_ ;
wire \u0_ps2_kb/_0071_ ;
wire \u0_ps2_kb/_0072_ ;
wire \u0_ps2_kb/_0073_ ;
wire \u0_ps2_kb/_0074_ ;
wire \u0_ps2_kb/_0075_ ;
wire \u0_ps2_kb/_0076_ ;
wire \u0_ps2_kb/_0077_ ;
wire \u0_ps2_kb/_0078_ ;
wire \u0_ps2_kb/_0079_ ;
wire \u0_ps2_kb/_0080_ ;
wire \u0_ps2_kb/_0081_ ;
wire \u0_ps2_kb/_0082_ ;
wire \u0_ps2_kb/_0083_ ;
wire \u0_ps2_kb/_0084_ ;
wire \u0_ps2_kb/_0085_ ;
wire \u0_ps2_kb/_0086_ ;
wire \u0_ps2_kb/_0087_ ;
wire \u0_ps2_kb/_0088_ ;
wire \u0_ps2_kb/_0089_ ;
wire \u0_ps2_kb/_0090_ ;
wire \u0_ps2_kb/_0091_ ;
wire \u0_ps2_kb/_0092_ ;
wire \u0_ps2_kb/_0093_ ;
wire \u0_ps2_kb/_0094_ ;
wire \u0_ps2_kb/_0095_ ;
wire \u0_ps2_kb/_0096_ ;
wire \u0_ps2_kb/_0097_ ;
wire \u0_ps2_kb/_0098_ ;
wire \u0_ps2_kb/_0099_ ;
wire \u0_ps2_kb/_0100_ ;
wire \u0_ps2_kb/_0101_ ;
wire \u0_ps2_kb/_0102_ ;
wire \u0_ps2_kb/_0103_ ;
wire \u0_ps2_kb/_0104_ ;
wire \u0_ps2_kb/_0105_ ;
wire \u0_ps2_kb/_0106_ ;
wire \u0_ps2_kb/_0107_ ;
wire \u0_ps2_kb/_0108_ ;
wire \u0_ps2_kb/_0109_ ;
wire \u0_ps2_kb/_0110_ ;
wire \u0_ps2_kb/_0111_ ;
wire \u0_ps2_kb/_0112_ ;
wire \u0_ps2_kb/_0113_ ;
wire \u0_ps2_kb/_0114_ ;
wire \u0_ps2_kb/_0115_ ;
wire \u0_ps2_kb/_0116_ ;
wire \u0_ps2_kb/_0117_ ;
wire \u0_ps2_kb/_0118_ ;
wire \u0_ps2_kb/_0119_ ;
wire \u0_ps2_kb/_0120_ ;
wire \u0_ps2_kb/_0121_ ;
wire \u0_ps2_kb/_0122_ ;
wire \u0_ps2_kb/_0123_ ;
wire \u0_ps2_kb/_0124_ ;
wire \u0_ps2_kb/_0125_ ;
wire \u0_ps2_kb/_0126_ ;
wire \u0_ps2_kb/_0127_ ;
wire \u0_ps2_kb/_0128_ ;
wire \u0_ps2_kb/_0129_ ;
wire \u0_ps2_kb/_0130_ ;
wire \u0_ps2_kb/_0131_ ;
wire \u0_ps2_kb/_0132_ ;
wire \u0_ps2_kb/_0133_ ;
wire \u0_ps2_kb/_0134_ ;
wire \u0_ps2_kb/_0135_ ;
wire \u0_ps2_kb/_0136_ ;
wire \u0_ps2_kb/_0137_ ;
wire \u0_ps2_kb/_0138_ ;
wire \u0_ps2_kb/_0139_ ;
wire \u0_ps2_kb/_0140_ ;
wire \u0_ps2_kb/_0141_ ;
wire \u0_ps2_kb/_0142_ ;
wire \u0_ps2_kb/_0143_ ;
wire \u0_ps2_kb/_0144_ ;
wire \u0_ps2_kb/_0145_ ;
wire \u0_ps2_kb/_0146_ ;
wire \u0_ps2_kb/_0147_ ;
wire \u0_ps2_kb/_0148_ ;
wire \u0_ps2_kb/_0149_ ;
wire \u0_ps2_kb/_0150_ ;
wire \u0_ps2_kb/_0151_ ;
wire \u0_ps2_kb/_0152_ ;
wire \u0_ps2_kb/_0153_ ;
wire \u0_ps2_kb/_0154_ ;
wire \u0_ps2_kb/_0155_ ;
wire \u0_ps2_kb/_0156_ ;
wire \u0_ps2_kb/_0157_ ;
wire \u0_ps2_kb/_0158_ ;
wire \u0_ps2_kb/_0159_ ;
wire \u0_ps2_kb/_0160_ ;
wire \u0_ps2_kb/_0161_ ;
wire \u0_ps2_kb/_0162_ ;
wire \u0_ps2_kb/_0163_ ;
wire \u0_ps2_kb/_0164_ ;
wire \u0_ps2_kb/_0165_ ;
wire \u0_ps2_kb/_0166_ ;
wire \u0_ps2_kb/_0167_ ;
wire \u0_ps2_kb/_0168_ ;
wire \u0_ps2_kb/_0169_ ;
wire \u0_ps2_kb/_0170_ ;
wire \u0_ps2_kb/_0171_ ;
wire \u0_ps2_kb/_0172_ ;
wire \u0_ps2_kb/_0173_ ;
wire \u0_ps2_kb/_0174_ ;
wire \u0_ps2_kb/_0175_ ;
wire \u0_ps2_kb/_0176_ ;
wire \u0_ps2_kb/_0177_ ;
wire \u0_ps2_kb/_0178_ ;
wire \u0_ps2_kb/_0179_ ;
wire \u0_ps2_kb/_0180_ ;
wire \u0_ps2_kb/_0181_ ;
wire \u0_ps2_kb/_0182_ ;
wire \u0_ps2_kb/_0183_ ;
wire \u0_ps2_kb/_0184_ ;
wire \u0_ps2_kb/_0185_ ;
wire \u0_ps2_kb/_0186_ ;
wire \u0_ps2_kb/_0187_ ;
wire \u0_ps2_kb/_0188_ ;
wire \u0_ps2_kb/_0189_ ;
wire \u0_ps2_kb/_0190_ ;
wire \u0_ps2_kb/_0191_ ;
wire \u0_ps2_kb/_0192_ ;
wire \u0_ps2_kb/_0193_ ;
wire \u0_ps2_kb/_0194_ ;
wire \u0_ps2_kb/_0195_ ;
wire \u0_ps2_kb/_0196_ ;
wire \u0_ps2_kb/_0197_ ;
wire \u0_ps2_kb/_0198_ ;
wire \u0_ps2_kb/_0199_ ;
wire \u0_ps2_kb/_0200_ ;
wire \u0_ps2_kb/_0201_ ;
wire \u0_ps2_kb/_0202_ ;
wire \u0_ps2_kb/_0203_ ;
wire \u0_ps2_kb/_0204_ ;
wire \u0_ps2_kb/_0205_ ;
wire \u0_ps2_kb/_0206_ ;
wire \u0_ps2_kb/_0207_ ;
wire \u0_ps2_kb/_0208_ ;
wire \u0_ps2_kb/_0209_ ;
wire \u0_ps2_kb/_0210_ ;
wire \u0_ps2_kb/_0211_ ;
wire \u0_ps2_kb/_0212_ ;
wire \u0_ps2_kb/_0213_ ;
wire \u0_ps2_kb/_0214_ ;
wire \u0_ps2_kb/_0215_ ;
wire \u0_ps2_kb/_0216_ ;
wire \u0_ps2_kb/_0217_ ;
wire \u0_ps2_kb/_0218_ ;
wire \u0_ps2_kb/_0219_ ;
wire \u0_ps2_kb/_0220_ ;
wire \u0_ps2_kb/_0221_ ;
wire \u0_ps2_kb/_0222_ ;
wire \u0_ps2_kb/_0223_ ;
wire \u0_ps2_kb/_0224_ ;
wire \u0_ps2_kb/_0225_ ;
wire \u0_ps2_kb/_0226_ ;
wire \u0_ps2_kb/_0227_ ;
wire \u0_ps2_kb/_0228_ ;
wire \u0_ps2_kb/_0229_ ;
wire \u0_ps2_kb/_0230_ ;
wire \u0_ps2_kb/_0231_ ;
wire \u0_ps2_kb/_0232_ ;
wire \u0_ps2_kb/_0233_ ;
wire \u0_ps2_kb/_0234_ ;
wire \u0_ps2_kb/_0235_ ;
wire \u0_ps2_kb/_0236_ ;
wire \u0_ps2_kb/_0237_ ;
wire \u0_ps2_kb/_0238_ ;
wire \u0_ps2_kb/_0239_ ;
wire \u0_ps2_kb/_0240_ ;
wire \u0_ps2_kb/_0241_ ;
wire \u0_ps2_kb/_0242_ ;
wire \u0_ps2_kb/_0243_ ;
wire \u0_ps2_kb/_0244_ ;
wire \u0_ps2_kb/_0245_ ;
wire \u0_ps2_kb/_0246_ ;
wire \u0_ps2_kb/_0247_ ;
wire \u0_ps2_kb/_0248_ ;
wire \u0_ps2_kb/_0249_ ;
wire \u0_ps2_kb/_0250_ ;
wire \u0_ps2_kb/_0251_ ;
wire \u0_ps2_kb/_0252_ ;
wire \u0_ps2_kb/_0253_ ;
wire \u0_ps2_kb/_0254_ ;
wire \u0_ps2_kb/_0255_ ;
wire \u0_ps2_kb/_0256_ ;
wire \u0_ps2_kb/_0257_ ;
wire \u0_ps2_kb/_0258_ ;
wire \u0_ps2_kb/_0259_ ;
wire \u0_ps2_kb/_0260_ ;
wire \u0_ps2_kb/_0261_ ;
wire \u0_ps2_kb/_0262_ ;
wire \u0_ps2_kb/_0263_ ;
wire \u0_ps2_kb/_0264_ ;
wire \u0_ps2_kb/_0265_ ;
wire \u0_ps2_kb/_0266_ ;
wire \u0_ps2_kb/_0267_ ;
wire \u0_ps2_kb/_0268_ ;
wire \u0_ps2_kb/_0269_ ;
wire \u0_ps2_kb/_0270_ ;
wire \u0_ps2_kb/_0271_ ;
wire \u0_ps2_kb/_0272_ ;
wire \u0_ps2_kb/_0273_ ;
wire \u0_ps2_kb/_0274_ ;
wire \u0_ps2_kb/_0275_ ;
wire \u0_ps2_kb/_0276_ ;
wire \u0_ps2_kb/_0277_ ;
wire \u0_ps2_kb/_0278_ ;
wire \u0_ps2_kb/_0279_ ;
wire \u0_ps2_kb/_0280_ ;
wire \u0_ps2_kb/_0281_ ;
wire \u0_ps2_kb/_0282_ ;
wire \u0_ps2_kb/_0283_ ;
wire \u0_ps2_kb/_0284_ ;
wire \u0_ps2_kb/_0285_ ;
wire \u0_ps2_kb/_0286_ ;
wire \u0_ps2_kb/_0287_ ;
wire \u0_ps2_kb/_0288_ ;
wire \u0_ps2_kb/_0289_ ;
wire \u0_ps2_kb/_0290_ ;
wire \u0_ps2_kb/_0291_ ;
wire \u0_ps2_kb/_0292_ ;
wire \u0_ps2_kb/_0293_ ;
wire \u0_ps2_kb/_0294_ ;
wire \u0_ps2_kb/_0295_ ;
wire \u0_ps2_kb/_0296_ ;
wire \u0_ps2_kb/_0297_ ;
wire \u0_ps2_kb/_0298_ ;
wire \u0_ps2_kb/_0299_ ;
wire \u0_ps2_kb/_0300_ ;
wire \u0_ps2_kb/_0301_ ;
wire \u0_ps2_kb/_0302_ ;
wire \u0_ps2_kb/_0303_ ;
wire \u0_ps2_kb/_0304_ ;
wire \u0_ps2_kb/_0305_ ;
wire \u0_ps2_kb/_0306_ ;
wire \u0_ps2_kb/_0307_ ;
wire \u0_ps2_kb/_0308_ ;
wire \u0_ps2_kb/_0309_ ;
wire \u0_ps2_kb/_0310_ ;
wire \u0_ps2_kb/_0311_ ;
wire \u0_ps2_kb/_0312_ ;
wire \u0_ps2_kb/_0313_ ;
wire \u0_ps2_kb/_0314_ ;
wire \u0_ps2_kb/_0315_ ;
wire \u0_ps2_kb/_0316_ ;
wire \u0_ps2_kb/_0317_ ;
wire \u0_ps2_kb/_0318_ ;
wire \u0_ps2_kb/_0319_ ;
wire \u0_ps2_kb/_0320_ ;
wire \u0_ps2_kb/_0321_ ;
wire \u0_ps2_kb/_0322_ ;
wire \u0_ps2_kb/_0323_ ;
wire \u0_ps2_kb/_0324_ ;
wire \u0_ps2_kb/_0325_ ;
wire \u0_ps2_kb/_0326_ ;
wire \u0_ps2_kb/_0327_ ;
wire \u0_ps2_kb/_0328_ ;
wire \u0_ps2_kb/_0329_ ;
wire \u0_ps2_kb/_0330_ ;
wire \u0_ps2_kb/_0331_ ;
wire \u0_ps2_kb/_0332_ ;
wire \u0_ps2_kb/_0333_ ;
wire \u0_ps2_kb/_0334_ ;
wire \u0_ps2_kb/_0335_ ;
wire \u0_ps2_kb/_0336_ ;
wire \u0_ps2_kb/_0337_ ;
wire \u0_ps2_kb/_0338_ ;
wire \u0_ps2_kb/_0339_ ;
wire \u0_ps2_kb/_0340_ ;
wire \u0_ps2_kb/_0341_ ;
wire \u0_ps2_kb/_0342_ ;
wire \u0_ps2_kb/_0343_ ;
wire \u0_ps2_kb/_0344_ ;
wire \u0_ps2_kb/_0345_ ;
wire \u0_ps2_kb/_0346_ ;
wire \u0_ps2_kb/_0347_ ;
wire \u0_ps2_kb/_0348_ ;
wire \u0_ps2_kb/_0349_ ;
wire \u0_ps2_kb/_0350_ ;
wire \u0_ps2_kb/_0351_ ;
wire \u0_ps2_kb/_0352_ ;
wire \u0_ps2_kb/_0353_ ;
wire \u0_ps2_kb/_0354_ ;
wire \u0_ps2_kb/_0355_ ;
wire \u0_ps2_kb/_0356_ ;
wire \u0_ps2_kb/_0357_ ;
wire \u0_ps2_kb/_0358_ ;
wire \u0_ps2_kb/_0359_ ;
wire \u0_ps2_kb/_0360_ ;
wire \u0_ps2_kb/_0361_ ;
wire \u0_ps2_kb/_0362_ ;
wire \u0_ps2_kb/_0363_ ;
wire \u0_ps2_kb/_0364_ ;
wire \u0_ps2_kb/_0365_ ;
wire \u0_ps2_kb/_0366_ ;
wire \u0_ps2_kb/_0367_ ;
wire \u0_ps2_kb/_0368_ ;
wire \u0_ps2_kb/_0369_ ;
wire \u0_ps2_kb/_0370_ ;
wire \u0_ps2_kb/_0371_ ;
wire \u0_ps2_kb/_0372_ ;
wire \u0_ps2_kb/_0373_ ;
wire \u0_ps2_kb/_0374_ ;
wire \u0_ps2_kb/_0375_ ;
wire \u0_ps2_kb/_0376_ ;
wire \u0_ps2_kb/_0377_ ;
wire \u0_ps2_kb/_0378_ ;
wire \u0_ps2_kb/_0379_ ;
wire \u0_ps2_kb/_0380_ ;
wire \u0_ps2_kb/_0381_ ;
wire \u0_ps2_kb/_0382_ ;
wire \u0_ps2_kb/_0383_ ;
wire \u0_ps2_kb/_0384_ ;
wire \u0_ps2_kb/_0385_ ;
wire \u0_ps2_kb/_0386_ ;
wire \u0_ps2_kb/_0387_ ;
wire \u0_ps2_kb/_0388_ ;
wire \u0_ps2_kb/_0389_ ;
wire \u0_ps2_kb/_0390_ ;
wire \u0_ps2_kb/_0391_ ;
wire \u0_ps2_kb/_0392_ ;
wire \u0_ps2_kb/_0393_ ;
wire \u0_ps2_kb/_0394_ ;
wire \u0_ps2_kb/_0395_ ;
wire \u0_ps2_kb/_0396_ ;
wire \u0_ps2_kb/_0397_ ;
wire \u0_ps2_kb/_0398_ ;
wire \u0_ps2_kb/_0399_ ;
wire \u0_ps2_kb/_0400_ ;
wire \u0_ps2_kb/_0401_ ;
wire \u0_ps2_kb/_0402_ ;
wire \u0_ps2_kb/_0403_ ;
wire \u0_ps2_kb/_0404_ ;
wire \u0_ps2_kb/_0405_ ;
wire \u0_ps2_kb/_0406_ ;
wire \u0_ps2_kb/_0407_ ;
wire \u0_ps2_kb/_0408_ ;
wire \u0_ps2_kb/_0409_ ;
wire \u0_ps2_kb/_0410_ ;
wire \u0_ps2_kb/_0411_ ;
wire \u0_ps2_kb/_0412_ ;
wire \u0_ps2_kb/_0413_ ;
wire \u0_ps2_kb/_0414_ ;
wire \u0_ps2_kb/_0415_ ;
wire \u0_ps2_kb/_0416_ ;
wire \u0_ps2_kb/_0417_ ;
wire \u0_ps2_kb/_0418_ ;
wire \u0_ps2_kb/_0419_ ;
wire \u0_ps2_kb/_0420_ ;
wire \u0_ps2_kb/_0421_ ;
wire \u0_ps2_kb/_0422_ ;
wire \u0_ps2_kb/_0423_ ;
wire \u0_ps2_kb/_0424_ ;
wire \u0_ps2_kb/_0425_ ;
wire \u0_ps2_kb/_0426_ ;
wire \u0_ps2_kb/_0427_ ;
wire \u0_ps2_kb/_0428_ ;
wire \u0_ps2_kb/_0429_ ;
wire \u0_ps2_kb/_0430_ ;
wire \u0_ps2_kb/_0431_ ;
wire \u0_ps2_kb/_0432_ ;
wire \u0_ps2_kb/_0433_ ;
wire \u0_ps2_kb/_0434_ ;
wire \u0_ps2_kb/_0435_ ;
wire \u0_ps2_kb/_0436_ ;
wire \u0_ps2_kb/_0437_ ;
wire \u0_ps2_kb/_0438_ ;
wire \u0_ps2_kb/_0439_ ;
wire \u0_ps2_kb/_0440_ ;
wire \u0_ps2_kb/_0441_ ;
wire \u0_ps2_kb/_0442_ ;
wire \u0_ps2_kb/_0443_ ;
wire \u0_ps2_kb/_0444_ ;
wire \u0_ps2_kb/_0445_ ;
wire \u0_ps2_kb/_0446_ ;
wire \u0_ps2_kb/_0447_ ;
wire \u0_ps2_kb/_0448_ ;
wire \u0_ps2_kb/_0449_ ;
wire \u0_ps2_kb/_0450_ ;
wire \u0_ps2_kb/_0451_ ;
wire \u0_ps2_kb/_0452_ ;
wire \u0_ps2_kb/_0453_ ;
wire \u0_ps2_kb/_0454_ ;
wire \u0_ps2_kb/_0455_ ;
wire \u0_ps2_kb/_0456_ ;
wire \u0_ps2_kb/_0457_ ;
wire \u0_ps2_kb/_0458_ ;
wire \u0_ps2_kb/_0459_ ;
wire \u0_ps2_kb/_0460_ ;
wire \u0_ps2_kb/_0461_ ;
wire \u0_ps2_kb/_0462_ ;
wire \u0_ps2_kb/_0463_ ;
wire \u0_ps2_kb/_0464_ ;
wire \u0_ps2_kb/_0465_ ;
wire \u0_ps2_kb/_0466_ ;
wire \u0_ps2_kb/_0467_ ;
wire \u0_ps2_kb/_0468_ ;
wire \u0_ps2_kb/_0469_ ;
wire \u0_ps2_kb/_0470_ ;
wire \u0_ps2_kb/_0471_ ;
wire \u0_ps2_kb/_0472_ ;
wire \u0_ps2_kb/_0473_ ;
wire \u0_ps2_kb/_0474_ ;
wire \u0_ps2_kb/_0475_ ;
wire \u0_ps2_kb/_0476_ ;
wire \u0_ps2_kb/_0477_ ;
wire \u0_ps2_kb/_0478_ ;
wire \u0_ps2_kb/_0479_ ;
wire \u0_ps2_kb/_0480_ ;
wire \u0_ps2_kb/_0481_ ;
wire \u0_ps2_kb/_0482_ ;
wire \u0_ps2_kb/_0483_ ;
wire \u0_ps2_kb/_0484_ ;
wire \u0_ps2_kb/_0485_ ;
wire \u0_ps2_kb/_0486_ ;
wire \u0_ps2_kb/_0487_ ;
wire \u0_ps2_kb/_0488_ ;
wire \u0_ps2_kb/_0489_ ;
wire \u0_ps2_kb/_0490_ ;
wire \u0_ps2_kb/_0491_ ;
wire \u0_ps2_kb/_0492_ ;
wire \u0_ps2_kb/_0493_ ;
wire \u0_ps2_kb/_0494_ ;
wire \u0_ps2_kb/_0495_ ;
wire \u0_ps2_kb/_0496_ ;
wire \u0_ps2_kb/_0497_ ;
wire \u0_ps2_kb/_0498_ ;
wire \u0_ps2_kb/_0499_ ;
wire \u0_ps2_kb/_0500_ ;
wire \u0_ps2_kb/_0501_ ;
wire \u0_ps2_kb/_0502_ ;
wire \u0_ps2_kb/_0503_ ;
wire \u0_ps2_kb/_0504_ ;
wire \u0_ps2_kb/_0505_ ;
wire \u0_ps2_kb/_0506_ ;
wire \u0_ps2_kb/_0507_ ;
wire \u0_ps2_kb/_0508_ ;
wire \u0_ps2_kb/_0509_ ;
wire \u0_ps2_kb/_0510_ ;
wire \u0_ps2_kb/_0511_ ;
wire \u0_ps2_kb/_0512_ ;
wire \u0_ps2_kb/_0513_ ;
wire \u0_ps2_kb/_0514_ ;
wire \u0_ps2_kb/_0515_ ;
wire \u0_ps2_kb/_0516_ ;
wire \u0_ps2_kb/_0517_ ;
wire \u0_ps2_kb/_0518_ ;
wire \u0_ps2_kb/_0519_ ;
wire \u0_ps2_kb/_0520_ ;
wire \u0_ps2_kb/_0521_ ;
wire \u0_ps2_kb/_0522_ ;
wire \u0_ps2_kb/_0523_ ;
wire \u0_ps2_kb/_0524_ ;
wire \u0_ps2_kb/_0525_ ;
wire \u0_ps2_kb/_0526_ ;
wire \u0_ps2_kb/_0527_ ;
wire \u0_ps2_kb/_0528_ ;
wire \u0_ps2_kb/_0529_ ;
wire \u0_ps2_kb/_0530_ ;
wire \u0_ps2_kb/_0531_ ;
wire \u0_ps2_kb/_0532_ ;
wire \u0_ps2_kb/_0533_ ;
wire \u0_ps2_kb/_0534_ ;
wire \u0_ps2_kb/_0535_ ;
wire \u0_ps2_kb/_0536_ ;
wire \u0_ps2_kb/_0537_ ;
wire \u0_ps2_kb/_0538_ ;
wire \u0_ps2_kb/_0539_ ;
wire \u0_ps2_kb/_0540_ ;
wire \u0_ps2_kb/_0541_ ;
wire \u0_ps2_kb/_0542_ ;
wire \u0_ps2_kb/_0543_ ;
wire \u0_ps2_kb/_0544_ ;
wire \u0_ps2_kb/_0545_ ;
wire \u0_ps2_kb/_0546_ ;
wire \u0_ps2_kb/_0547_ ;
wire \u0_ps2_kb/_0548_ ;
wire \u0_ps2_kb/_0549_ ;
wire \u0_ps2_kb/_0550_ ;
wire \u0_ps2_kb/_0551_ ;
wire \u0_ps2_kb/_0552_ ;
wire \u0_ps2_kb/_0553_ ;
wire \u0_ps2_kb/_0554_ ;
wire \u0_ps2_kb/_0555_ ;
wire \u0_ps2_kb/_0556_ ;
wire \u0_ps2_kb/_0557_ ;
wire \u0_ps2_kb/_0558_ ;
wire \u0_ps2_kb/_0559_ ;
wire \u0_ps2_kb/_0560_ ;
wire \u0_ps2_kb/_0561_ ;
wire \u0_ps2_kb/fifo[0][0] ;
wire \u0_ps2_kb/fifo[0][1] ;
wire \u0_ps2_kb/fifo[0][2] ;
wire \u0_ps2_kb/fifo[0][3] ;
wire \u0_ps2_kb/fifo[0][4] ;
wire \u0_ps2_kb/fifo[0][5] ;
wire \u0_ps2_kb/fifo[0][6] ;
wire \u0_ps2_kb/fifo[0][7] ;
wire \u0_ps2_kb/fifo[1][0] ;
wire \u0_ps2_kb/fifo[1][1] ;
wire \u0_ps2_kb/fifo[1][2] ;
wire \u0_ps2_kb/fifo[1][3] ;
wire \u0_ps2_kb/fifo[1][4] ;
wire \u0_ps2_kb/fifo[1][5] ;
wire \u0_ps2_kb/fifo[1][6] ;
wire \u0_ps2_kb/fifo[1][7] ;
wire \u0_ps2_kb/fifo[2][0] ;
wire \u0_ps2_kb/fifo[2][1] ;
wire \u0_ps2_kb/fifo[2][2] ;
wire \u0_ps2_kb/fifo[2][3] ;
wire \u0_ps2_kb/fifo[2][4] ;
wire \u0_ps2_kb/fifo[2][5] ;
wire \u0_ps2_kb/fifo[2][6] ;
wire \u0_ps2_kb/fifo[2][7] ;
wire \u0_ps2_kb/fifo[3][0] ;
wire \u0_ps2_kb/fifo[3][1] ;
wire \u0_ps2_kb/fifo[3][2] ;
wire \u0_ps2_kb/fifo[3][3] ;
wire \u0_ps2_kb/fifo[3][4] ;
wire \u0_ps2_kb/fifo[3][5] ;
wire \u0_ps2_kb/fifo[3][6] ;
wire \u0_ps2_kb/fifo[3][7] ;
wire \u0_ps2_kb/fifo[4][0] ;
wire \u0_ps2_kb/fifo[4][1] ;
wire \u0_ps2_kb/fifo[4][2] ;
wire \u0_ps2_kb/fifo[4][3] ;
wire \u0_ps2_kb/fifo[4][4] ;
wire \u0_ps2_kb/fifo[4][5] ;
wire \u0_ps2_kb/fifo[4][6] ;
wire \u0_ps2_kb/fifo[4][7] ;
wire \u0_ps2_kb/fifo[5][0] ;
wire \u0_ps2_kb/fifo[5][1] ;
wire \u0_ps2_kb/fifo[5][2] ;
wire \u0_ps2_kb/fifo[5][3] ;
wire \u0_ps2_kb/fifo[5][4] ;
wire \u0_ps2_kb/fifo[5][5] ;
wire \u0_ps2_kb/fifo[5][6] ;
wire \u0_ps2_kb/fifo[5][7] ;
wire \u0_ps2_kb/fifo[6][0] ;
wire \u0_ps2_kb/fifo[6][1] ;
wire \u0_ps2_kb/fifo[6][2] ;
wire \u0_ps2_kb/fifo[6][3] ;
wire \u0_ps2_kb/fifo[6][4] ;
wire \u0_ps2_kb/fifo[6][5] ;
wire \u0_ps2_kb/fifo[6][6] ;
wire \u0_ps2_kb/fifo[6][7] ;
wire \u0_ps2_kb/fifo[7][0] ;
wire \u0_ps2_kb/fifo[7][1] ;
wire \u0_ps2_kb/fifo[7][2] ;
wire \u0_ps2_kb/fifo[7][3] ;
wire \u0_ps2_kb/fifo[7][4] ;
wire \u0_ps2_kb/fifo[7][5] ;
wire \u0_ps2_kb/fifo[7][6] ;
wire \u0_ps2_kb/fifo[7][7] ;
wire \u1_ps2_dsh/_000_ ;
wire \u1_ps2_dsh/_001_ ;
wire \u1_ps2_dsh/_002_ ;
wire \u1_ps2_dsh/_003_ ;
wire \u1_ps2_dsh/_004_ ;
wire \u1_ps2_dsh/_005_ ;
wire \u1_ps2_dsh/_006_ ;
wire \u1_ps2_dsh/_007_ ;
wire \u1_ps2_dsh/_008_ ;
wire \u1_ps2_dsh/_009_ ;
wire \u1_ps2_dsh/_010_ ;
wire \u1_ps2_dsh/_011_ ;
wire \u1_ps2_dsh/_012_ ;
wire \u1_ps2_dsh/_013_ ;
wire \u1_ps2_dsh/_014_ ;
wire \u1_ps2_dsh/_015_ ;
wire \u1_ps2_dsh/_016_ ;
wire \u1_ps2_dsh/_017_ ;
wire \u1_ps2_dsh/_018_ ;
wire \u1_ps2_dsh/_019_ ;
wire \u1_ps2_dsh/_020_ ;
wire \u1_ps2_dsh/_021_ ;
wire \u1_ps2_dsh/_022_ ;
wire \u1_ps2_dsh/_023_ ;
wire \u1_ps2_dsh/_024_ ;
wire \u1_ps2_dsh/_025_ ;
wire \u1_ps2_dsh/_026_ ;
wire \u1_ps2_dsh/_027_ ;
wire \u1_ps2_dsh/_028_ ;
wire \u1_ps2_dsh/_029_ ;
wire \u1_ps2_dsh/_030_ ;
wire \u1_ps2_dsh/_031_ ;
wire \u1_ps2_dsh/_032_ ;
wire \u1_ps2_dsh/_033_ ;
wire \u1_ps2_dsh/_034_ ;
wire \u1_ps2_dsh/_035_ ;
wire \u1_ps2_dsh/_036_ ;
wire \u1_ps2_dsh/_037_ ;
wire \u1_ps2_dsh/_038_ ;
wire \u1_ps2_dsh/_039_ ;
wire \u1_ps2_dsh/_040_ ;
wire \u1_ps2_dsh/_041_ ;
wire \u1_ps2_dsh/_042_ ;
wire \u1_ps2_dsh/_043_ ;
wire \u1_ps2_dsh/_044_ ;
wire \u1_ps2_dsh/_045_ ;
wire \u1_ps2_dsh/_046_ ;
wire \u1_ps2_dsh/_047_ ;
wire \u1_ps2_dsh/_048_ ;
wire \u1_ps2_dsh/_049_ ;
wire \u1_ps2_dsh/_050_ ;
wire \u1_ps2_dsh/_051_ ;
wire \u2_ps2_cer/_000_ ;
wire \u2_ps2_cer/_001_ ;
wire \u2_ps2_cer/_002_ ;
wire \u2_ps2_cer/_003_ ;
wire \u2_ps2_cer/_004_ ;
wire \u2_ps2_cer/_005_ ;
wire \u2_ps2_cer/_006_ ;
wire \u2_ps2_cer/_007_ ;
wire \u2_ps2_cer/_008_ ;
wire \u2_ps2_cer/_009_ ;
wire \u2_ps2_cer/_010_ ;
wire \u2_ps2_cer/_011_ ;
wire \u2_ps2_cer/_012_ ;
wire \u2_ps2_cer/_013_ ;
wire \u2_ps2_cer/_014_ ;
wire \u2_ps2_cer/_015_ ;
wire \u2_ps2_cer/_016_ ;
wire \u2_ps2_cer/_017_ ;
wire \u2_ps2_cer/_018_ ;
wire \u2_ps2_cer/_019_ ;
wire \u2_ps2_cer/_020_ ;
wire \u2_ps2_cer/_021_ ;
wire \u2_ps2_cer/_022_ ;
wire \u2_ps2_cer/_023_ ;
wire \u2_ps2_cer/_024_ ;
wire \u2_ps2_cer/_025_ ;
wire \u2_ps2_cer/_026_ ;
wire \u2_ps2_cer/_027_ ;
wire \u2_ps2_cer/_028_ ;
wire \u2_ps2_cer/_029_ ;
wire \u2_ps2_cer/_030_ ;
wire \u2_ps2_cer/_031_ ;
wire \u2_ps2_cer/_032_ ;
wire \u2_ps2_cer/_033_ ;
wire \u2_ps2_cer/_034_ ;
wire \u2_ps2_cer/_035_ ;
wire \u2_ps2_cer/_036_ ;
wire \u2_ps2_cer/_037_ ;
wire \u2_ps2_cer/_038_ ;
wire \u2_ps2_cer/_039_ ;
wire \u2_ps2_cer/_040_ ;
wire \u2_ps2_cer/_041_ ;
wire \u2_ps2_cer/_042_ ;
wire \u2_ps2_cer/_043_ ;
wire \u2_ps2_cer/_044_ ;
wire \u2_ps2_cer/_045_ ;
wire \u2_ps2_cer/_046_ ;
wire \u2_ps2_cer/_047_ ;
wire \u2_ps2_cer/_048_ ;
wire \u2_ps2_cer/_049_ ;
wire \u2_ps2_cer/_050_ ;
wire \u2_ps2_cer/_051_ ;
wire \u2_ps2_cer/_052_ ;
wire \u2_ps2_cer/_053_ ;
wire \u2_ps2_cer/_054_ ;
wire \u2_ps2_cer/_055_ ;
wire \u2_ps2_cer/_056_ ;
wire \u2_ps2_cer/_057_ ;
wire \u2_ps2_cer/_058_ ;
wire \u2_ps2_cer/_059_ ;
wire \u2_ps2_cer/_060_ ;
wire \u2_ps2_cer/_061_ ;
wire \u2_ps2_cer/_062_ ;
wire \u2_ps2_cer/_063_ ;
wire \u2_ps2_cer/_064_ ;
wire \u2_ps2_cer/_065_ ;
wire \u2_ps2_cer/_066_ ;
wire \u2_ps2_cer/counted ;
wire \u3_seg_h_0/_00_ ;
wire \u3_seg_h_0/_01_ ;
wire \u3_seg_h_0/_02_ ;
wire \u3_seg_h_0/_03_ ;
wire \u3_seg_h_0/_04_ ;
wire \u3_seg_h_0/_05_ ;
wire \u3_seg_h_0/_06_ ;
wire \u3_seg_h_0/_07_ ;
wire \u3_seg_h_0/_08_ ;
wire \u3_seg_h_0/_09_ ;
wire \u3_seg_h_0/_10_ ;
wire \u3_seg_h_0/_11_ ;
wire \u3_seg_h_0/_12_ ;
wire \u3_seg_h_0/_13_ ;
wire \u3_seg_h_0/_14_ ;
wire \u3_seg_h_0/_15_ ;
wire \u3_seg_h_0/_16_ ;
wire \u3_seg_h_0/_17_ ;
wire \u3_seg_h_0/_18_ ;
wire \u3_seg_h_0/_19_ ;
wire \u3_seg_h_0/_20_ ;
wire \u3_seg_h_0/_21_ ;
wire \u3_seg_h_0/_22_ ;
wire \u3_seg_h_0/_23_ ;
wire \u3_seg_h_0/_24_ ;
wire \u3_seg_h_0/_25_ ;
wire \u3_seg_h_0/_26_ ;
wire \u3_seg_h_0/_27_ ;
wire \u3_seg_h_0/_28_ ;
wire \u3_seg_h_0/_29_ ;
wire \u3_seg_h_0/_30_ ;
wire \u3_seg_h_0/_31_ ;
wire \u3_seg_h_0/_32_ ;
wire \u3_seg_h_0/_33_ ;
wire \u3_seg_h_0/_34_ ;
wire \u3_seg_h_0/_35_ ;
wire \u3_seg_h_0/_36_ ;
wire \u3_seg_h_0/_37_ ;
wire \u3_seg_h_0/_38_ ;
wire \u3_seg_h_0/_39_ ;
wire \u3_seg_h_0/_40_ ;
wire \u3_seg_h_0/_41_ ;
wire \u3_seg_h_0/_42_ ;
wire \u4_seg_h_1/_00_ ;
wire \u4_seg_h_1/_01_ ;
wire \u4_seg_h_1/_02_ ;
wire \u4_seg_h_1/_03_ ;
wire \u4_seg_h_1/_04_ ;
wire \u4_seg_h_1/_05_ ;
wire \u4_seg_h_1/_06_ ;
wire \u4_seg_h_1/_07_ ;
wire \u4_seg_h_1/_08_ ;
wire \u4_seg_h_1/_09_ ;
wire \u4_seg_h_1/_10_ ;
wire \u4_seg_h_1/_11_ ;
wire \u4_seg_h_1/_12_ ;
wire \u4_seg_h_1/_13_ ;
wire \u4_seg_h_1/_14_ ;
wire \u4_seg_h_1/_15_ ;
wire \u4_seg_h_1/_16_ ;
wire \u4_seg_h_1/_17_ ;
wire \u4_seg_h_1/_18_ ;
wire \u4_seg_h_1/_19_ ;
wire \u4_seg_h_1/_20_ ;
wire \u4_seg_h_1/_21_ ;
wire \u4_seg_h_1/_22_ ;
wire \u4_seg_h_1/_23_ ;
wire \u4_seg_h_1/_24_ ;
wire \u4_seg_h_1/_25_ ;
wire \u4_seg_h_1/_26_ ;
wire \u4_seg_h_1/_27_ ;
wire \u4_seg_h_1/_28_ ;
wire \u4_seg_h_1/_29_ ;
wire \u4_seg_h_1/_30_ ;
wire \u4_seg_h_1/_31_ ;
wire \u4_seg_h_1/_32_ ;
wire \u4_seg_h_1/_33_ ;
wire \u4_seg_h_1/_34_ ;
wire \u4_seg_h_1/_35_ ;
wire \u4_seg_h_1/_36_ ;
wire \u4_seg_h_1/_37_ ;
wire \u4_seg_h_1/_38_ ;
wire \u4_seg_h_1/_39_ ;
wire \u4_seg_h_1/_40_ ;
wire \u4_seg_h_1/_41_ ;
wire \u4_seg_h_1/_42_ ;
wire \u5_seg_h_2/_00_ ;
wire \u5_seg_h_2/_01_ ;
wire \u5_seg_h_2/_02_ ;
wire \u5_seg_h_2/_03_ ;
wire \u5_seg_h_2/_04_ ;
wire \u5_seg_h_2/_05_ ;
wire \u5_seg_h_2/_06_ ;
wire \u5_seg_h_2/_07_ ;
wire \u5_seg_h_2/_08_ ;
wire \u5_seg_h_2/_09_ ;
wire \u5_seg_h_2/_10_ ;
wire \u5_seg_h_2/_11_ ;
wire \u5_seg_h_2/_12_ ;
wire \u5_seg_h_2/_13_ ;
wire \u5_seg_h_2/_14_ ;
wire \u5_seg_h_2/_15_ ;
wire \u5_seg_h_2/_16_ ;
wire \u5_seg_h_2/_17_ ;
wire \u5_seg_h_2/_18_ ;
wire \u5_seg_h_2/_19_ ;
wire \u5_seg_h_2/_20_ ;
wire \u5_seg_h_2/_21_ ;
wire \u5_seg_h_2/_22_ ;
wire \u5_seg_h_2/_23_ ;
wire \u5_seg_h_2/_24_ ;
wire \u5_seg_h_2/_25_ ;
wire \u5_seg_h_2/_26_ ;
wire \u5_seg_h_2/_27_ ;
wire \u5_seg_h_2/_28_ ;
wire \u5_seg_h_2/_29_ ;
wire \u5_seg_h_2/_30_ ;
wire \u5_seg_h_2/_31_ ;
wire \u5_seg_h_2/_32_ ;
wire \u5_seg_h_2/_33_ ;
wire \u5_seg_h_2/_34_ ;
wire \u5_seg_h_2/_35_ ;
wire \u5_seg_h_2/_36_ ;
wire \u5_seg_h_2/_37_ ;
wire \u5_seg_h_2/_38_ ;
wire \u5_seg_h_2/_39_ ;
wire \u5_seg_h_2/_40_ ;
wire \u5_seg_h_2/_41_ ;
wire \u5_seg_h_2/_42_ ;
wire \u6_seg_h_3/_00_ ;
wire \u6_seg_h_3/_01_ ;
wire \u6_seg_h_3/_02_ ;
wire \u6_seg_h_3/_03_ ;
wire \u6_seg_h_3/_04_ ;
wire \u6_seg_h_3/_05_ ;
wire \u6_seg_h_3/_06_ ;
wire \u6_seg_h_3/_07_ ;
wire \u6_seg_h_3/_08_ ;
wire \u6_seg_h_3/_09_ ;
wire \u6_seg_h_3/_10_ ;
wire \u6_seg_h_3/_11_ ;
wire \u6_seg_h_3/_12_ ;
wire \u6_seg_h_3/_13_ ;
wire \u6_seg_h_3/_14_ ;
wire \u6_seg_h_3/_15_ ;
wire \u6_seg_h_3/_16_ ;
wire \u6_seg_h_3/_17_ ;
wire \u6_seg_h_3/_18_ ;
wire \u6_seg_h_3/_19_ ;
wire \u6_seg_h_3/_20_ ;
wire \u6_seg_h_3/_21_ ;
wire \u6_seg_h_3/_22_ ;
wire \u6_seg_h_3/_23_ ;
wire \u6_seg_h_3/_24_ ;
wire \u6_seg_h_3/_25_ ;
wire \u6_seg_h_3/_26_ ;
wire \u6_seg_h_3/_27_ ;
wire \u6_seg_h_3/_28_ ;
wire \u6_seg_h_3/_29_ ;
wire \u6_seg_h_3/_30_ ;
wire \u6_seg_h_3/_31_ ;
wire \u6_seg_h_3/_32_ ;
wire \u6_seg_h_3/_33_ ;
wire \u6_seg_h_3/_34_ ;
wire \u6_seg_h_3/_35_ ;
wire \u6_seg_h_3/_36_ ;
wire \u6_seg_h_3/_37_ ;
wire \u6_seg_h_3/_38_ ;
wire \u6_seg_h_3/_39_ ;
wire \u6_seg_h_3/_40_ ;
wire \u6_seg_h_3/_41_ ;
wire \u6_seg_h_3/_42_ ;
wire \u7_seg_h_4/_00_ ;
wire \u7_seg_h_4/_01_ ;
wire \u7_seg_h_4/_02_ ;
wire \u7_seg_h_4/_03_ ;
wire \u7_seg_h_4/_04_ ;
wire \u7_seg_h_4/_05_ ;
wire \u7_seg_h_4/_06_ ;
wire \u7_seg_h_4/_07_ ;
wire \u7_seg_h_4/_08_ ;
wire \u7_seg_h_4/_09_ ;
wire \u7_seg_h_4/_10_ ;
wire \u7_seg_h_4/_11_ ;
wire \u7_seg_h_4/_12_ ;
wire \u7_seg_h_4/_13_ ;
wire \u7_seg_h_4/_14_ ;
wire \u7_seg_h_4/_15_ ;
wire \u7_seg_h_4/_16_ ;
wire \u7_seg_h_4/_17_ ;
wire \u7_seg_h_4/_18_ ;
wire \u7_seg_h_4/_19_ ;
wire \u7_seg_h_4/_20_ ;
wire \u7_seg_h_4/_21_ ;
wire \u7_seg_h_4/_22_ ;
wire \u7_seg_h_4/_23_ ;
wire \u7_seg_h_4/_24_ ;
wire \u7_seg_h_4/_25_ ;
wire \u7_seg_h_4/_26_ ;
wire \u7_seg_h_4/_27_ ;
wire \u7_seg_h_4/_28_ ;
wire \u7_seg_h_4/_29_ ;
wire \u7_seg_h_4/_30_ ;
wire \u7_seg_h_4/_31_ ;
wire \u7_seg_h_4/_32_ ;
wire \u7_seg_h_4/_33_ ;
wire \u7_seg_h_4/_34_ ;
wire \u7_seg_h_4/_35_ ;
wire \u7_seg_h_4/_36_ ;
wire \u7_seg_h_4/_37_ ;
wire \u7_seg_h_4/_38_ ;
wire \u7_seg_h_4/_39_ ;
wire \u7_seg_h_4/_40_ ;
wire \u7_seg_h_4/_41_ ;
wire \u7_seg_h_4/_42_ ;
wire \u8_seg_h_5/_00_ ;
wire \u8_seg_h_5/_01_ ;
wire \u8_seg_h_5/_02_ ;
wire \u8_seg_h_5/_03_ ;
wire \u8_seg_h_5/_04_ ;
wire \u8_seg_h_5/_05_ ;
wire \u8_seg_h_5/_06_ ;
wire \u8_seg_h_5/_07_ ;
wire \u8_seg_h_5/_08_ ;
wire \u8_seg_h_5/_09_ ;
wire \u8_seg_h_5/_10_ ;
wire \u8_seg_h_5/_11_ ;
wire \u8_seg_h_5/_12_ ;
wire \u8_seg_h_5/_13_ ;
wire \u8_seg_h_5/_14_ ;
wire \u8_seg_h_5/_15_ ;
wire \u8_seg_h_5/_16_ ;
wire \u8_seg_h_5/_17_ ;
wire \u8_seg_h_5/_18_ ;
wire \u8_seg_h_5/_19_ ;
wire \u8_seg_h_5/_20_ ;
wire \u8_seg_h_5/_21_ ;
wire \u8_seg_h_5/_22_ ;
wire \u8_seg_h_5/_23_ ;
wire \u8_seg_h_5/_24_ ;
wire \u8_seg_h_5/_25_ ;
wire \u8_seg_h_5/_26_ ;
wire \u8_seg_h_5/_27_ ;
wire \u8_seg_h_5/_28_ ;
wire \u8_seg_h_5/_29_ ;
wire \u8_seg_h_5/_30_ ;
wire \u8_seg_h_5/_31_ ;
wire \u8_seg_h_5/_32_ ;
wire \u8_seg_h_5/_33_ ;
wire \u8_seg_h_5/_34_ ;
wire \u8_seg_h_5/_35_ ;
wire \u8_seg_h_5/_36_ ;
wire \u8_seg_h_5/_37_ ;
wire \u8_seg_h_5/_38_ ;
wire \u8_seg_h_5/_39_ ;
wire \u8_seg_h_5/_40_ ;
wire \u8_seg_h_5/_41_ ;
wire \u8_seg_h_5/_42_ ;
wire clk ;
wire clrn ;
wire ps2_data ;
wire overflow ;
wire ps2_clk ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire \ascii[0] ;
wire \ascii[1] ;
wire \ascii[2] ;
wire \ascii[3] ;
wire \ascii[4] ;
wire \ascii[5] ;
wire \ascii[6] ;
wire \ascii[7] ;
wire \data[0] ;
wire \data[1] ;
wire \data[2] ;
wire \data[3] ;
wire \data[4] ;
wire \data[5] ;
wire \data[6] ;
wire \data[7] ;
wire \data_d1[0] ;
wire \data_d1[1] ;
wire \data_d1[2] ;
wire \data_d1[3] ;
wire \data_d1[4] ;
wire \data_d1[5] ;
wire \data_d1[6] ;
wire \data_d1[7] ;
wire \high_tens[0] ;
wire \high_tens[1] ;
wire \high_tens[2] ;
wire \high_tens[3] ;
wire \high_units[0] ;
wire \high_units[1] ;
wire \high_units[2] ;
wire \high_units[3] ;
wire \key_ascii_display[0] ;
wire \key_ascii_display[1] ;
wire \key_ascii_display[2] ;
wire \key_ascii_display[3] ;
wire \key_ascii_display[4] ;
wire \key_ascii_display[5] ;
wire \key_ascii_display[6] ;
wire \key_ascii_display[7] ;
wire \key_scan_display[0] ;
wire \key_scan_display[1] ;
wire \key_scan_display[2] ;
wire \key_scan_display[3] ;
wire \key_scan_display[4] ;
wire \key_scan_display[5] ;
wire \key_scan_display[6] ;
wire \key_scan_display[7] ;
wire \u0_ps2_kb/buffer[0] ;
wire \u0_ps2_kb/buffer[1] ;
wire \u0_ps2_kb/buffer[2] ;
wire \u0_ps2_kb/buffer[3] ;
wire \u0_ps2_kb/buffer[4] ;
wire \u0_ps2_kb/buffer[5] ;
wire \u0_ps2_kb/buffer[6] ;
wire \u0_ps2_kb/buffer[7] ;
wire \u0_ps2_kb/buffer[8] ;
wire \u0_ps2_kb/buffer[9] ;
wire \u0_ps2_kb/count[0] ;
wire \u0_ps2_kb/count[1] ;
wire \u0_ps2_kb/count[2] ;
wire \u0_ps2_kb/count[3] ;
wire \u0_ps2_kb/ps2_clk_sync[0] ;
wire \u0_ps2_kb/ps2_clk_sync[1] ;
wire \u0_ps2_kb/ps2_clk_sync[2] ;
wire \u0_ps2_kb/r_ptr[0] ;
wire \u0_ps2_kb/r_ptr[1] ;
wire \u0_ps2_kb/r_ptr[2] ;
wire \u0_ps2_kb/w_ptr[0] ;
wire \u0_ps2_kb/w_ptr[1] ;
wire \u0_ps2_kb/w_ptr[2] ;
wire \u1_ps2_dsh/ascii_result[0] ;
wire \u1_ps2_dsh/ascii_result[1] ;
wire \u1_ps2_dsh/ascii_result[2] ;
wire \u1_ps2_dsh/ascii_result[3] ;
wire \u1_ps2_dsh/ascii_result[4] ;
wire \u1_ps2_dsh/ascii_result[5] ;
wire \u1_ps2_dsh/ascii_result[6] ;
wire \u1_ps2_dsh/ascii_result[7] ;
wire \seg_out_2[0] ;
wire \seg_out_2[1] ;
wire \seg_out_2[2] ;
wire \seg_out_2[3] ;
wire \seg_out_2[4] ;
wire \seg_out_2[5] ;
wire \seg_out_2[6] ;
wire \seg_out_2[7] ;
wire \seg_out_3[0] ;
wire \seg_out_3[1] ;
wire \seg_out_3[2] ;
wire \seg_out_3[3] ;
wire \seg_out_3[4] ;
wire \seg_out_3[5] ;
wire \seg_out_3[6] ;
wire \seg_out_3[7] ;
wire \seg_out_0[0] ;
wire \seg_out_0[1] ;
wire \seg_out_0[2] ;
wire \seg_out_0[3] ;
wire \seg_out_0[4] ;
wire \seg_out_0[5] ;
wire \seg_out_0[6] ;
wire \seg_out_0[7] ;
wire \seg_out_1[0] ;
wire \seg_out_1[1] ;
wire \seg_out_1[2] ;
wire \seg_out_1[3] ;
wire \seg_out_1[4] ;
wire \seg_out_1[5] ;
wire \seg_out_1[6] ;
wire \seg_out_1[7] ;
wire \seg_out_4[0] ;
wire \seg_out_4[1] ;
wire \seg_out_4[2] ;
wire \seg_out_4[3] ;
wire \seg_out_4[4] ;
wire \seg_out_4[5] ;
wire \seg_out_4[6] ;
wire \seg_out_4[7] ;
wire \seg_out_5[0] ;
wire \seg_out_5[1] ;
wire \seg_out_5[2] ;
wire \seg_out_5[3] ;
wire \seg_out_5[4] ;
wire \seg_out_5[5] ;
wire \seg_out_5[6] ;
wire \seg_out_5[7] ;

assign seg_out_2[0] = \seg_out_2[0] ;
assign seg_out_2[1] = \seg_out_2[1] ;
assign seg_out_2[2] = \seg_out_2[2] ;
assign seg_out_2[3] = \seg_out_2[3] ;
assign seg_out_2[4] = \seg_out_2[4] ;
assign seg_out_2[5] = \seg_out_2[5] ;
assign seg_out_2[6] = \seg_out_2[6] ;
assign seg_out_2[7] = \seg_out_2[7] ;
assign seg_out_3[0] = \seg_out_3[0] ;
assign seg_out_3[1] = \seg_out_3[1] ;
assign seg_out_3[2] = \seg_out_3[2] ;
assign seg_out_3[3] = \seg_out_3[3] ;
assign seg_out_3[4] = \seg_out_3[4] ;
assign seg_out_3[5] = \seg_out_3[5] ;
assign seg_out_3[6] = \seg_out_3[6] ;
assign seg_out_3[7] = \seg_out_3[7] ;
assign seg_out_0[0] = \seg_out_0[0] ;
assign seg_out_0[1] = \seg_out_0[1] ;
assign seg_out_0[2] = \seg_out_0[2] ;
assign seg_out_0[3] = \seg_out_0[3] ;
assign seg_out_0[4] = \seg_out_0[4] ;
assign seg_out_0[5] = \seg_out_0[5] ;
assign seg_out_0[6] = \seg_out_0[6] ;
assign seg_out_0[7] = \seg_out_0[7] ;
assign seg_out_1[0] = \seg_out_1[0] ;
assign seg_out_1[1] = \seg_out_1[1] ;
assign seg_out_1[2] = \seg_out_1[2] ;
assign seg_out_1[3] = \seg_out_1[3] ;
assign seg_out_1[4] = \seg_out_1[4] ;
assign seg_out_1[5] = \seg_out_1[5] ;
assign seg_out_1[6] = \seg_out_1[6] ;
assign seg_out_1[7] = \seg_out_1[7] ;
assign seg_out_4[0] = \seg_out_4[0] ;
assign seg_out_4[1] = \seg_out_4[1] ;
assign seg_out_4[2] = \seg_out_4[2] ;
assign seg_out_4[3] = \seg_out_4[3] ;
assign seg_out_4[4] = \seg_out_4[4] ;
assign seg_out_4[5] = \seg_out_4[5] ;
assign seg_out_4[6] = \seg_out_4[6] ;
assign seg_out_4[7] = \seg_out_4[7] ;
assign seg_out_5[0] = \seg_out_5[0] ;
assign seg_out_5[1] = \seg_out_5[1] ;
assign seg_out_5[2] = \seg_out_5[2] ;
assign seg_out_5[3] = \seg_out_5[3] ;
assign seg_out_5[4] = \seg_out_5[4] ;
assign seg_out_5[5] = \seg_out_5[5] ;
assign seg_out_5[6] = \seg_out_5[6] ;
assign seg_out_5[7] = \seg_out_5[7] ;

INV_X32 _133_ ( .A(_103_ ), .ZN(_098_ ) );
NOR3_X1 _134_ ( .A1(_098_ ), .A2(_104_ ), .A3(_087_ ), .ZN(_053_ ) );
NOR2_X4 _135_ ( .A1(_098_ ), .A2(_104_ ), .ZN(_099_ ) );
BUF_X4 _136_ ( .A(_099_ ), .Z(_100_ ) );
MUX2_X1 _137_ ( .A(_070_ ), .B(_062_ ), .S(_100_ ), .Z(_027_ ) );
MUX2_X1 _138_ ( .A(_071_ ), .B(_063_ ), .S(_100_ ), .Z(_028_ ) );
MUX2_X1 _139_ ( .A(_072_ ), .B(_064_ ), .S(_100_ ), .Z(_029_ ) );
MUX2_X1 _140_ ( .A(_073_ ), .B(_065_ ), .S(_100_ ), .Z(_030_ ) );
MUX2_X1 _141_ ( .A(_074_ ), .B(_066_ ), .S(_100_ ), .Z(_031_ ) );
MUX2_X1 _142_ ( .A(_075_ ), .B(_067_ ), .S(_100_ ), .Z(_032_ ) );
MUX2_X1 _143_ ( .A(_076_ ), .B(_068_ ), .S(_100_ ), .Z(_033_ ) );
MUX2_X1 _144_ ( .A(_077_ ), .B(_069_ ), .S(_100_ ), .Z(_034_ ) );
MUX2_X1 _145_ ( .A(_079_ ), .B(_054_ ), .S(_100_ ), .Z(_036_ ) );
BUF_X4 _146_ ( .A(_099_ ), .Z(_101_ ) );
MUX2_X1 _147_ ( .A(_080_ ), .B(_055_ ), .S(_101_ ), .Z(_037_ ) );
MUX2_X1 _148_ ( .A(_081_ ), .B(_056_ ), .S(_101_ ), .Z(_038_ ) );
MUX2_X1 _149_ ( .A(_082_ ), .B(_057_ ), .S(_101_ ), .Z(_039_ ) );
MUX2_X1 _150_ ( .A(_083_ ), .B(_058_ ), .S(_101_ ), .Z(_040_ ) );
MUX2_X1 _151_ ( .A(_084_ ), .B(_059_ ), .S(_101_ ), .Z(_041_ ) );
MUX2_X1 _152_ ( .A(_085_ ), .B(_060_ ), .S(_101_ ), .Z(_042_ ) );
MUX2_X1 _153_ ( .A(_086_ ), .B(_061_ ), .S(_101_ ), .Z(_043_ ) );
MUX2_X1 _154_ ( .A(_088_ ), .B(_062_ ), .S(_101_ ), .Z(_044_ ) );
MUX2_X1 _155_ ( .A(_089_ ), .B(_063_ ), .S(_101_ ), .Z(_045_ ) );
MUX2_X1 _156_ ( .A(_090_ ), .B(_064_ ), .S(_101_ ), .Z(_046_ ) );
MUX2_X1 _157_ ( .A(_091_ ), .B(_065_ ), .S(_099_ ), .Z(_047_ ) );
MUX2_X1 _158_ ( .A(_092_ ), .B(_066_ ), .S(_099_ ), .Z(_048_ ) );
MUX2_X1 _159_ ( .A(_093_ ), .B(_067_ ), .S(_099_ ), .Z(_049_ ) );
MUX2_X1 _160_ ( .A(_094_ ), .B(_068_ ), .S(_099_ ), .Z(_050_ ) );
MUX2_X1 _161_ ( .A(_095_ ), .B(_069_ ), .S(_099_ ), .Z(_051_ ) );
INV_X1 _162_ ( .A(_102_ ), .ZN(_096_ ) );
AOI21_X1 _163_ ( .A(_100_ ), .B1(_087_ ), .B2(_096_ ), .ZN(_052_ ) );
INV_X1 _164_ ( .A(_078_ ), .ZN(_097_ ) );
OAI22_X1 _165_ ( .A1(_098_ ), .A2(_104_ ), .B1(_097_ ), .B2(_087_ ), .ZN(_035_ ) );
LOGIC1_X1 _166_ ( .Z(_132_ ) );
BUF_X1 _167_ ( .A(ready ), .Z(_103_ ) );
BUF_X1 _168_ ( .A(ready_d1 ), .Z(_104_ ) );
BUF_X1 _169_ ( .A(key_release ), .Z(_087_ ) );
BUF_X1 _170_ ( .A(_053_ ), .Z(_026_ ) );
BUF_X1 _171_ ( .A(\data[0] ), .Z(_062_ ) );
BUF_X1 _172_ ( .A(\data_d1[0] ), .Z(_070_ ) );
BUF_X1 _173_ ( .A(_027_ ), .Z(_000_ ) );
BUF_X1 _174_ ( .A(\data[1] ), .Z(_063_ ) );
BUF_X1 _175_ ( .A(\data_d1[1] ), .Z(_071_ ) );
BUF_X1 _176_ ( .A(_028_ ), .Z(_001_ ) );
BUF_X1 _177_ ( .A(\data[2] ), .Z(_064_ ) );
BUF_X1 _178_ ( .A(\data_d1[2] ), .Z(_072_ ) );
BUF_X1 _179_ ( .A(_029_ ), .Z(_002_ ) );
BUF_X1 _180_ ( .A(\data[3] ), .Z(_065_ ) );
BUF_X1 _181_ ( .A(\data_d1[3] ), .Z(_073_ ) );
BUF_X1 _182_ ( .A(_030_ ), .Z(_003_ ) );
BUF_X1 _183_ ( .A(\data[4] ), .Z(_066_ ) );
BUF_X1 _184_ ( .A(\data_d1[4] ), .Z(_074_ ) );
BUF_X1 _185_ ( .A(_031_ ), .Z(_004_ ) );
BUF_X1 _186_ ( .A(\data[5] ), .Z(_067_ ) );
BUF_X1 _187_ ( .A(\data_d1[5] ), .Z(_075_ ) );
BUF_X1 _188_ ( .A(_032_ ), .Z(_005_ ) );
BUF_X1 _189_ ( .A(\data[6] ), .Z(_068_ ) );
BUF_X1 _190_ ( .A(\data_d1[6] ), .Z(_076_ ) );
BUF_X1 _191_ ( .A(_033_ ), .Z(_006_ ) );
BUF_X1 _192_ ( .A(\data[7] ), .Z(_069_ ) );
BUF_X1 _193_ ( .A(\data_d1[7] ), .Z(_077_ ) );
BUF_X1 _194_ ( .A(_034_ ), .Z(_007_ ) );
BUF_X1 _195_ ( .A(\ascii[0] ), .Z(_054_ ) );
BUF_X1 _196_ ( .A(\key_ascii_display[0] ), .Z(_079_ ) );
BUF_X1 _197_ ( .A(_036_ ), .Z(_009_ ) );
BUF_X1 _198_ ( .A(\ascii[1] ), .Z(_055_ ) );
BUF_X1 _199_ ( .A(\key_ascii_display[1] ), .Z(_080_ ) );
BUF_X1 _200_ ( .A(_037_ ), .Z(_010_ ) );
BUF_X1 _201_ ( .A(\ascii[2] ), .Z(_056_ ) );
BUF_X1 _202_ ( .A(\key_ascii_display[2] ), .Z(_081_ ) );
BUF_X1 _203_ ( .A(_038_ ), .Z(_011_ ) );
BUF_X1 _204_ ( .A(\ascii[3] ), .Z(_057_ ) );
BUF_X1 _205_ ( .A(\key_ascii_display[3] ), .Z(_082_ ) );
BUF_X1 _206_ ( .A(_039_ ), .Z(_012_ ) );
BUF_X1 _207_ ( .A(\ascii[4] ), .Z(_058_ ) );
BUF_X1 _208_ ( .A(\key_ascii_display[4] ), .Z(_083_ ) );
BUF_X1 _209_ ( .A(_040_ ), .Z(_013_ ) );
BUF_X1 _210_ ( .A(\ascii[5] ), .Z(_059_ ) );
BUF_X1 _211_ ( .A(\key_ascii_display[5] ), .Z(_084_ ) );
BUF_X1 _212_ ( .A(_041_ ), .Z(_014_ ) );
BUF_X1 _213_ ( .A(\ascii[6] ), .Z(_060_ ) );
BUF_X1 _214_ ( .A(\key_ascii_display[6] ), .Z(_085_ ) );
BUF_X1 _215_ ( .A(_042_ ), .Z(_015_ ) );
BUF_X1 _216_ ( .A(\ascii[7] ), .Z(_061_ ) );
BUF_X1 _217_ ( .A(\key_ascii_display[7] ), .Z(_086_ ) );
BUF_X1 _218_ ( .A(_043_ ), .Z(_016_ ) );
BUF_X1 _219_ ( .A(\key_scan_display[0] ), .Z(_088_ ) );
BUF_X1 _220_ ( .A(_044_ ), .Z(_017_ ) );
BUF_X1 _221_ ( .A(\key_scan_display[1] ), .Z(_089_ ) );
BUF_X1 _222_ ( .A(_045_ ), .Z(_018_ ) );
BUF_X1 _223_ ( .A(\key_scan_display[2] ), .Z(_090_ ) );
BUF_X1 _224_ ( .A(_046_ ), .Z(_019_ ) );
BUF_X1 _225_ ( .A(\key_scan_display[3] ), .Z(_091_ ) );
BUF_X1 _226_ ( .A(_047_ ), .Z(_020_ ) );
BUF_X1 _227_ ( .A(\key_scan_display[4] ), .Z(_092_ ) );
BUF_X1 _228_ ( .A(_048_ ), .Z(_021_ ) );
BUF_X1 _229_ ( .A(\key_scan_display[5] ), .Z(_093_ ) );
BUF_X1 _230_ ( .A(_049_ ), .Z(_022_ ) );
BUF_X1 _231_ ( .A(\key_scan_display[6] ), .Z(_094_ ) );
BUF_X1 _232_ ( .A(_050_ ), .Z(_023_ ) );
BUF_X1 _233_ ( .A(\key_scan_display[7] ), .Z(_095_ ) );
BUF_X1 _234_ ( .A(_051_ ), .Z(_024_ ) );
BUF_X1 _235_ ( .A(nextdata_n ), .Z(_102_ ) );
BUF_X1 _236_ ( .A(_052_ ), .Z(_025_ ) );
BUF_X1 _237_ ( .A(en ), .Z(_078_ ) );
BUF_X1 _238_ ( .A(_035_ ), .Z(_008_ ) );
DFFS_X1 _239_ ( .D(_025_ ), .SN(fanout_net_2 ), .CK(clk ), .Q(nextdata_n ), .QN(_105_ ) );
DFFR_X1 _240_ ( .D(_000_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[0] ), .QN(_106_ ) );
DFFR_X1 _241_ ( .D(_001_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[1] ), .QN(_107_ ) );
DFFR_X1 _242_ ( .D(_002_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[2] ), .QN(_108_ ) );
DFFR_X1 _243_ ( .D(_003_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[3] ), .QN(_109_ ) );
DFFR_X1 _244_ ( .D(_004_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[4] ), .QN(_110_ ) );
DFFR_X1 _245_ ( .D(_005_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[5] ), .QN(_111_ ) );
DFFR_X1 _246_ ( .D(_006_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[6] ), .QN(_112_ ) );
DFFR_X1 _247_ ( .D(_007_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\data_d1[7] ), .QN(_113_ ) );
DFFR_X1 _248_ ( .D(_017_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[0] ), .QN(_114_ ) );
DFFR_X1 _249_ ( .D(_018_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[1] ), .QN(_115_ ) );
DFFR_X1 _250_ ( .D(_019_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[2] ), .QN(_116_ ) );
DFFR_X1 _251_ ( .D(_020_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[3] ), .QN(_117_ ) );
DFFR_X1 _252_ ( .D(_021_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[4] ), .QN(_118_ ) );
DFFR_X1 _253_ ( .D(_022_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[5] ), .QN(_119_ ) );
DFFR_X1 _254_ ( .D(_023_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[6] ), .QN(_120_ ) );
DFFR_X1 _255_ ( .D(_024_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_scan_display[7] ), .QN(_121_ ) );
DFFR_X1 _256_ ( .D(_009_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[0] ), .QN(_122_ ) );
DFFR_X1 _257_ ( .D(_010_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[1] ), .QN(_123_ ) );
DFFR_X1 _258_ ( .D(_011_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[2] ), .QN(_124_ ) );
DFFR_X1 _259_ ( .D(_012_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[3] ), .QN(_125_ ) );
DFFR_X1 _260_ ( .D(_013_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[4] ), .QN(_126_ ) );
DFFR_X1 _261_ ( .D(_014_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[5] ), .QN(_127_ ) );
DFFR_X1 _262_ ( .D(_015_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[6] ), .QN(_128_ ) );
DFFR_X1 _263_ ( .D(_016_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\key_ascii_display[7] ), .QN(_129_ ) );
DFFR_X1 _264_ ( .D(_008_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(en ), .QN(_130_ ) );
DFFR_X1 _265_ ( .D(ready ), .RN(fanout_net_2 ), .CK(clk ), .Q(ready_d1 ), .QN(_131_ ) );
INV_X1 \u0_ps2_kb/_0562_ ( .A(\u0_ps2_kb/_0474_ ), .ZN(\u0_ps2_kb/_0279_ ) );
NOR2_X1 \u0_ps2_kb/_0563_ ( .A1(\u0_ps2_kb/_0279_ ), .A2(\u0_ps2_kb/_0473_ ), .ZN(\u0_ps2_kb/_0280_ ) );
INV_X1 \u0_ps2_kb/_0564_ ( .A(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0281_ ) );
NOR2_X1 \u0_ps2_kb/_0565_ ( .A1(\u0_ps2_kb/_0281_ ), .A2(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0282_ ) );
AND2_X1 \u0_ps2_kb/_0566_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0282_ ), .ZN(\u0_ps2_kb/_0283_ ) );
INV_X1 \u0_ps2_kb/_0567_ ( .A(\u0_ps2_kb/_0206_ ), .ZN(\u0_ps2_kb/_0284_ ) );
NAND2_X1 \u0_ps2_kb/_0568_ ( .A1(\u0_ps2_kb/_0284_ ), .A2(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0285_ ) );
INV_X1 \u0_ps2_kb/_0569_ ( .A(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0286_ ) );
NOR2_X1 \u0_ps2_kb/_0570_ ( .A1(\u0_ps2_kb/_0285_ ), .A2(\u0_ps2_kb/_0286_ ), .ZN(\u0_ps2_kb/_0287_ ) );
NAND2_X1 \u0_ps2_kb/_0571_ ( .A1(\u0_ps2_kb/_0283_ ), .A2(\u0_ps2_kb/_0287_ ), .ZN(\u0_ps2_kb/_0288_ ) );
MUX2_X1 \u0_ps2_kb/_0572_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0288_ ), .Z(\u0_ps2_kb/_0102_ ) );
AND2_X1 \u0_ps2_kb/_0573_ ( .A1(\u0_ps2_kb/_0203_ ), .A2(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0289_ ) );
AND2_X1 \u0_ps2_kb/_0574_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0289_ ), .ZN(\u0_ps2_kb/_0290_ ) );
NAND2_X1 \u0_ps2_kb/_0575_ ( .A1(\u0_ps2_kb/_0290_ ), .A2(\u0_ps2_kb/_0287_ ), .ZN(\u0_ps2_kb/_0291_ ) );
MUX2_X1 \u0_ps2_kb/_0576_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0291_ ), .Z(\u0_ps2_kb/_0103_ ) );
INV_X1 \u0_ps2_kb/_0577_ ( .A(\u0_ps2_kb/_0475_ ), .ZN(\u0_ps2_kb/_0292_ ) );
XOR2_X2 \u0_ps2_kb/_0578_ ( .A(\u0_ps2_kb/_0196_ ), .B(\u0_ps2_kb/_0195_ ), .Z(\u0_ps2_kb/_0293_ ) );
XNOR2_X2 \u0_ps2_kb/_0579_ ( .A(\u0_ps2_kb/_0198_ ), .B(\u0_ps2_kb/_0199_ ), .ZN(\u0_ps2_kb/_0294_ ) );
XNOR2_X2 \u0_ps2_kb/_0580_ ( .A(\u0_ps2_kb/_0293_ ), .B(\u0_ps2_kb/_0294_ ), .ZN(\u0_ps2_kb/_0295_ ) );
XNOR2_X1 \u0_ps2_kb/_0581_ ( .A(\u0_ps2_kb/_0194_ ), .B(\u0_ps2_kb/_0193_ ), .ZN(\u0_ps2_kb/_0296_ ) );
XNOR2_X2 \u0_ps2_kb/_0582_ ( .A(\u0_ps2_kb/_0197_ ), .B(\u0_ps2_kb/_0200_ ), .ZN(\u0_ps2_kb/_0297_ ) );
XNOR2_X1 \u0_ps2_kb/_0583_ ( .A(\u0_ps2_kb/_0296_ ), .B(\u0_ps2_kb/_0297_ ), .ZN(\u0_ps2_kb/_0298_ ) );
XNOR2_X2 \u0_ps2_kb/_0584_ ( .A(\u0_ps2_kb/_0295_ ), .B(\u0_ps2_kb/_0298_ ), .ZN(\u0_ps2_kb/_0299_ ) );
AOI211_X2 \u0_ps2_kb/_0585_ ( .A(\u0_ps2_kb/_0292_ ), .B(\u0_ps2_kb/_0192_ ), .C1(\u0_ps2_kb/_0299_ ), .C2(\u0_ps2_kb/_0201_ ), .ZN(\u0_ps2_kb/_0300_ ) );
OR2_X1 \u0_ps2_kb/_0586_ ( .A1(\u0_ps2_kb/_0299_ ), .A2(\u0_ps2_kb/_0201_ ), .ZN(\u0_ps2_kb/_0301_ ) );
AND2_X2 \u0_ps2_kb/_0587_ ( .A1(\u0_ps2_kb/_0300_ ), .A2(\u0_ps2_kb/_0301_ ), .ZN(\u0_ps2_kb/_0302_ ) );
NOR2_X1 \u0_ps2_kb/_0588_ ( .A1(\u0_ps2_kb/_0284_ ), .A2(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0303_ ) );
AND2_X1 \u0_ps2_kb/_0589_ ( .A1(\u0_ps2_kb/_0282_ ), .A2(\u0_ps2_kb/_0303_ ), .ZN(\u0_ps2_kb/_0304_ ) );
AND2_X1 \u0_ps2_kb/_0590_ ( .A1(\u0_ps2_kb/_0304_ ), .A2(\u0_ps2_kb/_0280_ ), .ZN(\u0_ps2_kb/_0305_ ) );
AND2_X4 \u0_ps2_kb/_0591_ ( .A1(\u0_ps2_kb/_0302_ ), .A2(\u0_ps2_kb/_0305_ ), .ZN(\u0_ps2_kb/_0306_ ) );
NAND2_X4 \u0_ps2_kb/_0592_ ( .A1(\u0_ps2_kb/_0306_ ), .A2(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0307_ ) );
BUF_X16 \u0_ps2_kb/_0593_ ( .A(\u0_ps2_kb/_0307_ ), .Z(\u0_ps2_kb/_0308_ ) );
BUF_X8 \u0_ps2_kb/_0594_ ( .A(\u0_ps2_kb/_0308_ ), .Z(\u0_ps2_kb/_0309_ ) );
INV_X1 \u0_ps2_kb/_0595_ ( .A(\u0_ps2_kb/_0482_ ), .ZN(\u0_ps2_kb/_0310_ ) );
NAND3_X1 \u0_ps2_kb/_0596_ ( .A1(\u0_ps2_kb/_0310_ ), .A2(\u0_ps2_kb/_0481_ ), .A3(\u0_ps2_kb/_0480_ ), .ZN(\u0_ps2_kb/_0311_ ) );
NOR3_X1 \u0_ps2_kb/_0597_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0193_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0312_ ) );
INV_X1 \u0_ps2_kb/_0598_ ( .A(\u0_ps2_kb/_0239_ ), .ZN(\u0_ps2_kb/_0313_ ) );
OR2_X4 \u0_ps2_kb/_0599_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0314_ ) );
AOI21_X1 \u0_ps2_kb/_0600_ ( .A(\u0_ps2_kb/_0312_ ), .B1(\u0_ps2_kb/_0313_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0142_ ) );
NOR3_X1 \u0_ps2_kb/_0601_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0194_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0315_ ) );
INV_X1 \u0_ps2_kb/_0602_ ( .A(\u0_ps2_kb/_0240_ ), .ZN(\u0_ps2_kb/_0316_ ) );
AOI21_X1 \u0_ps2_kb/_0603_ ( .A(\u0_ps2_kb/_0315_ ), .B1(\u0_ps2_kb/_0316_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0143_ ) );
NOR3_X1 \u0_ps2_kb/_0604_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0195_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0317_ ) );
INV_X1 \u0_ps2_kb/_0605_ ( .A(\u0_ps2_kb/_0241_ ), .ZN(\u0_ps2_kb/_0318_ ) );
AOI21_X1 \u0_ps2_kb/_0606_ ( .A(\u0_ps2_kb/_0317_ ), .B1(\u0_ps2_kb/_0318_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0144_ ) );
NOR3_X1 \u0_ps2_kb/_0607_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0196_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0319_ ) );
INV_X1 \u0_ps2_kb/_0608_ ( .A(\u0_ps2_kb/_0242_ ), .ZN(\u0_ps2_kb/_0320_ ) );
AOI21_X1 \u0_ps2_kb/_0609_ ( .A(\u0_ps2_kb/_0319_ ), .B1(\u0_ps2_kb/_0320_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0145_ ) );
NOR2_X4 \u0_ps2_kb/_0610_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0321_ ) );
MUX2_X1 \u0_ps2_kb/_0611_ ( .A(\u0_ps2_kb/_0243_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0321_ ), .Z(\u0_ps2_kb/_0146_ ) );
MUX2_X1 \u0_ps2_kb/_0612_ ( .A(\u0_ps2_kb/_0244_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0321_ ), .Z(\u0_ps2_kb/_0147_ ) );
NOR3_X1 \u0_ps2_kb/_0613_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0199_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0322_ ) );
INV_X1 \u0_ps2_kb/_0614_ ( .A(\u0_ps2_kb/_0245_ ), .ZN(\u0_ps2_kb/_0323_ ) );
AOI21_X1 \u0_ps2_kb/_0615_ ( .A(\u0_ps2_kb/_0322_ ), .B1(\u0_ps2_kb/_0323_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0148_ ) );
NOR3_X1 \u0_ps2_kb/_0616_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0200_ ), .A3(\u0_ps2_kb/_0311_ ), .ZN(\u0_ps2_kb/_0324_ ) );
INV_X1 \u0_ps2_kb/_0617_ ( .A(\u0_ps2_kb/_0246_ ), .ZN(\u0_ps2_kb/_0325_ ) );
AOI21_X1 \u0_ps2_kb/_0618_ ( .A(\u0_ps2_kb/_0324_ ), .B1(\u0_ps2_kb/_0325_ ), .B2(\u0_ps2_kb/_0314_ ), .ZN(\u0_ps2_kb/_0149_ ) );
INV_X1 \u0_ps2_kb/_0619_ ( .A(\u0_ps2_kb/_0481_ ), .ZN(\u0_ps2_kb/_0326_ ) );
INV_X1 \u0_ps2_kb/_0620_ ( .A(\u0_ps2_kb/_0480_ ), .ZN(\u0_ps2_kb/_0327_ ) );
NAND3_X1 \u0_ps2_kb/_0621_ ( .A1(\u0_ps2_kb/_0326_ ), .A2(\u0_ps2_kb/_0327_ ), .A3(\u0_ps2_kb/_0482_ ), .ZN(\u0_ps2_kb/_0328_ ) );
NOR2_X4 \u0_ps2_kb/_0622_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0328_ ), .ZN(\u0_ps2_kb/_0329_ ) );
MUX2_X1 \u0_ps2_kb/_0623_ ( .A(\u0_ps2_kb/_0247_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0150_ ) );
MUX2_X1 \u0_ps2_kb/_0624_ ( .A(\u0_ps2_kb/_0248_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0151_ ) );
MUX2_X1 \u0_ps2_kb/_0625_ ( .A(\u0_ps2_kb/_0249_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0152_ ) );
MUX2_X1 \u0_ps2_kb/_0626_ ( .A(\u0_ps2_kb/_0250_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0153_ ) );
MUX2_X1 \u0_ps2_kb/_0627_ ( .A(\u0_ps2_kb/_0251_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0154_ ) );
MUX2_X1 \u0_ps2_kb/_0628_ ( .A(\u0_ps2_kb/_0252_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0155_ ) );
MUX2_X1 \u0_ps2_kb/_0629_ ( .A(\u0_ps2_kb/_0253_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0156_ ) );
MUX2_X1 \u0_ps2_kb/_0630_ ( .A(\u0_ps2_kb/_0254_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0329_ ), .Z(\u0_ps2_kb/_0157_ ) );
NAND3_X1 \u0_ps2_kb/_0631_ ( .A1(\u0_ps2_kb/_0310_ ), .A2(\u0_ps2_kb/_0326_ ), .A3(\u0_ps2_kb/_0327_ ), .ZN(\u0_ps2_kb/_0330_ ) );
NOR2_X2 \u0_ps2_kb/_0632_ ( .A1(\u0_ps2_kb/_0307_ ), .A2(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0331_ ) );
MUX2_X1 \u0_ps2_kb/_0633_ ( .A(\u0_ps2_kb/_0215_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0118_ ) );
MUX2_X1 \u0_ps2_kb/_0634_ ( .A(\u0_ps2_kb/_0216_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0119_ ) );
MUX2_X1 \u0_ps2_kb/_0635_ ( .A(\u0_ps2_kb/_0217_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0120_ ) );
MUX2_X1 \u0_ps2_kb/_0636_ ( .A(\u0_ps2_kb/_0218_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0121_ ) );
NOR3_X1 \u0_ps2_kb/_0637_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0197_ ), .A3(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0332_ ) );
INV_X1 \u0_ps2_kb/_0638_ ( .A(\u0_ps2_kb/_0219_ ), .ZN(\u0_ps2_kb/_0333_ ) );
OR2_X2 \u0_ps2_kb/_0639_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0334_ ) );
AOI21_X1 \u0_ps2_kb/_0640_ ( .A(\u0_ps2_kb/_0332_ ), .B1(\u0_ps2_kb/_0333_ ), .B2(\u0_ps2_kb/_0334_ ), .ZN(\u0_ps2_kb/_0122_ ) );
NOR3_X1 \u0_ps2_kb/_0641_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0198_ ), .A3(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0335_ ) );
INV_X1 \u0_ps2_kb/_0642_ ( .A(\u0_ps2_kb/_0220_ ), .ZN(\u0_ps2_kb/_0336_ ) );
AOI21_X1 \u0_ps2_kb/_0643_ ( .A(\u0_ps2_kb/_0335_ ), .B1(\u0_ps2_kb/_0336_ ), .B2(\u0_ps2_kb/_0334_ ), .ZN(\u0_ps2_kb/_0123_ ) );
MUX2_X1 \u0_ps2_kb/_0644_ ( .A(\u0_ps2_kb/_0221_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0331_ ), .Z(\u0_ps2_kb/_0124_ ) );
NOR3_X1 \u0_ps2_kb/_0645_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0200_ ), .A3(\u0_ps2_kb/_0330_ ), .ZN(\u0_ps2_kb/_0337_ ) );
INV_X1 \u0_ps2_kb/_0646_ ( .A(\u0_ps2_kb/_0222_ ), .ZN(\u0_ps2_kb/_0338_ ) );
AOI21_X1 \u0_ps2_kb/_0647_ ( .A(\u0_ps2_kb/_0337_ ), .B1(\u0_ps2_kb/_0338_ ), .B2(\u0_ps2_kb/_0334_ ), .ZN(\u0_ps2_kb/_0125_ ) );
INV_X1 \u0_ps2_kb/_0648_ ( .A(\u0_ps2_kb/_0477_ ), .ZN(\u0_ps2_kb/_0339_ ) );
BUF_X2 \u0_ps2_kb/_0649_ ( .A(\u0_ps2_kb/_0339_ ), .Z(\u0_ps2_kb/_0340_ ) );
NOR2_X1 \u0_ps2_kb/_0650_ ( .A1(fanout_net_1 ), .A2(\u0_ps2_kb/_0231_ ), .ZN(\u0_ps2_kb/_0341_ ) );
AOI211_X4 \u0_ps2_kb/_0651_ ( .A(\u0_ps2_kb/_0340_ ), .B(\u0_ps2_kb/_0341_ ), .C1(\u0_ps2_kb/_0313_ ), .C2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0342_ ) );
MUX2_X1 \u0_ps2_kb/_0652_ ( .A(\u0_ps2_kb/_0215_ ), .B(\u0_ps2_kb/_0223_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0343_ ) );
AOI211_X4 \u0_ps2_kb/_0653_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0342_ ), .C1(\u0_ps2_kb/_0340_ ), .C2(\u0_ps2_kb/_0343_ ), .ZN(\u0_ps2_kb/_0344_ ) );
MUX2_X1 \u0_ps2_kb/_0654_ ( .A(\u0_ps2_kb/_0255_ ), .B(\u0_ps2_kb/_0271_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0345_ ) );
AND2_X1 \u0_ps2_kb/_0655_ ( .A1(\u0_ps2_kb/_0345_ ), .A2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0346_ ) );
INV_X1 \u0_ps2_kb/_0656_ ( .A(fanout_net_1 ), .ZN(\u0_ps2_kb/_0347_ ) );
MUX2_X1 \u0_ps2_kb/_0657_ ( .A(\u0_ps2_kb/_0247_ ), .B(\u0_ps2_kb/_0263_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0348_ ) );
AOI21_X1 \u0_ps2_kb/_0658_ ( .A(\u0_ps2_kb/_0346_ ), .B1(\u0_ps2_kb/_0347_ ), .B2(\u0_ps2_kb/_0348_ ), .ZN(\u0_ps2_kb/_0349_ ) );
AOI21_X1 \u0_ps2_kb/_0659_ ( .A(\u0_ps2_kb/_0344_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0349_ ), .ZN(\u0_ps2_kb/_0207_ ) );
NOR2_X1 \u0_ps2_kb/_0660_ ( .A1(fanout_net_1 ), .A2(\u0_ps2_kb/_0232_ ), .ZN(\u0_ps2_kb/_0350_ ) );
AOI211_X4 \u0_ps2_kb/_0661_ ( .A(\u0_ps2_kb/_0340_ ), .B(\u0_ps2_kb/_0350_ ), .C1(\u0_ps2_kb/_0316_ ), .C2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0351_ ) );
MUX2_X1 \u0_ps2_kb/_0662_ ( .A(\u0_ps2_kb/_0216_ ), .B(\u0_ps2_kb/_0224_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0352_ ) );
AOI211_X4 \u0_ps2_kb/_0663_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0351_ ), .C1(\u0_ps2_kb/_0340_ ), .C2(\u0_ps2_kb/_0352_ ), .ZN(\u0_ps2_kb/_0353_ ) );
MUX2_X1 \u0_ps2_kb/_0664_ ( .A(\u0_ps2_kb/_0248_ ), .B(\u0_ps2_kb/_0264_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0354_ ) );
AND2_X1 \u0_ps2_kb/_0665_ ( .A1(\u0_ps2_kb/_0354_ ), .A2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0355_ ) );
MUX2_X1 \u0_ps2_kb/_0666_ ( .A(\u0_ps2_kb/_0256_ ), .B(\u0_ps2_kb/_0272_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0356_ ) );
AOI21_X1 \u0_ps2_kb/_0667_ ( .A(\u0_ps2_kb/_0355_ ), .B1(fanout_net_1 ), .B2(\u0_ps2_kb/_0356_ ), .ZN(\u0_ps2_kb/_0357_ ) );
AOI21_X1 \u0_ps2_kb/_0668_ ( .A(\u0_ps2_kb/_0353_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0357_ ), .ZN(\u0_ps2_kb/_0208_ ) );
NOR2_X1 \u0_ps2_kb/_0669_ ( .A1(fanout_net_1 ), .A2(\u0_ps2_kb/_0233_ ), .ZN(\u0_ps2_kb/_0358_ ) );
AOI211_X4 \u0_ps2_kb/_0670_ ( .A(\u0_ps2_kb/_0340_ ), .B(\u0_ps2_kb/_0358_ ), .C1(\u0_ps2_kb/_0318_ ), .C2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0359_ ) );
MUX2_X1 \u0_ps2_kb/_0671_ ( .A(\u0_ps2_kb/_0217_ ), .B(\u0_ps2_kb/_0225_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0360_ ) );
AOI211_X4 \u0_ps2_kb/_0672_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0359_ ), .C1(\u0_ps2_kb/_0340_ ), .C2(\u0_ps2_kb/_0360_ ), .ZN(\u0_ps2_kb/_0361_ ) );
MUX2_X1 \u0_ps2_kb/_0673_ ( .A(\u0_ps2_kb/_0249_ ), .B(\u0_ps2_kb/_0265_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0362_ ) );
AND2_X1 \u0_ps2_kb/_0674_ ( .A1(\u0_ps2_kb/_0362_ ), .A2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0363_ ) );
MUX2_X1 \u0_ps2_kb/_0675_ ( .A(\u0_ps2_kb/_0257_ ), .B(\u0_ps2_kb/_0273_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0364_ ) );
AOI21_X1 \u0_ps2_kb/_0676_ ( .A(\u0_ps2_kb/_0363_ ), .B1(fanout_net_1 ), .B2(\u0_ps2_kb/_0364_ ), .ZN(\u0_ps2_kb/_0365_ ) );
AOI21_X1 \u0_ps2_kb/_0677_ ( .A(\u0_ps2_kb/_0361_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0365_ ), .ZN(\u0_ps2_kb/_0209_ ) );
NOR2_X1 \u0_ps2_kb/_0678_ ( .A1(fanout_net_1 ), .A2(\u0_ps2_kb/_0234_ ), .ZN(\u0_ps2_kb/_0366_ ) );
AOI211_X4 \u0_ps2_kb/_0679_ ( .A(\u0_ps2_kb/_0340_ ), .B(\u0_ps2_kb/_0366_ ), .C1(\u0_ps2_kb/_0320_ ), .C2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0367_ ) );
MUX2_X1 \u0_ps2_kb/_0680_ ( .A(\u0_ps2_kb/_0218_ ), .B(\u0_ps2_kb/_0226_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0368_ ) );
AOI211_X4 \u0_ps2_kb/_0681_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0367_ ), .C1(\u0_ps2_kb/_0340_ ), .C2(\u0_ps2_kb/_0368_ ), .ZN(\u0_ps2_kb/_0369_ ) );
MUX2_X1 \u0_ps2_kb/_0682_ ( .A(\u0_ps2_kb/_0250_ ), .B(\u0_ps2_kb/_0258_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0370_ ) );
AND2_X1 \u0_ps2_kb/_0683_ ( .A1(\u0_ps2_kb/_0370_ ), .A2(\u0_ps2_kb/_0340_ ), .ZN(\u0_ps2_kb/_0371_ ) );
MUX2_X1 \u0_ps2_kb/_0684_ ( .A(\u0_ps2_kb/_0266_ ), .B(\u0_ps2_kb/_0274_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0372_ ) );
AOI21_X1 \u0_ps2_kb/_0685_ ( .A(\u0_ps2_kb/_0371_ ), .B1(\u0_ps2_kb/_0477_ ), .B2(\u0_ps2_kb/_0372_ ), .ZN(\u0_ps2_kb/_0373_ ) );
AOI21_X1 \u0_ps2_kb/_0686_ ( .A(\u0_ps2_kb/_0369_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0373_ ), .ZN(\u0_ps2_kb/_0210_ ) );
NOR2_X1 \u0_ps2_kb/_0687_ ( .A1(\u0_ps2_kb/_0347_ ), .A2(\u0_ps2_kb/_0227_ ), .ZN(\u0_ps2_kb/_0374_ ) );
AOI211_X4 \u0_ps2_kb/_0688_ ( .A(\u0_ps2_kb/_0477_ ), .B(\u0_ps2_kb/_0374_ ), .C1(\u0_ps2_kb/_0333_ ), .C2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0375_ ) );
MUX2_X1 \u0_ps2_kb/_0689_ ( .A(\u0_ps2_kb/_0235_ ), .B(\u0_ps2_kb/_0243_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0376_ ) );
AOI211_X4 \u0_ps2_kb/_0690_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0375_ ), .C1(\u0_ps2_kb/_0477_ ), .C2(\u0_ps2_kb/_0376_ ), .ZN(\u0_ps2_kb/_0377_ ) );
MUX2_X1 \u0_ps2_kb/_0691_ ( .A(\u0_ps2_kb/_0251_ ), .B(\u0_ps2_kb/_0267_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0378_ ) );
AND2_X1 \u0_ps2_kb/_0692_ ( .A1(\u0_ps2_kb/_0378_ ), .A2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0379_ ) );
MUX2_X1 \u0_ps2_kb/_0693_ ( .A(\u0_ps2_kb/_0259_ ), .B(\u0_ps2_kb/_0275_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0380_ ) );
AOI21_X1 \u0_ps2_kb/_0694_ ( .A(\u0_ps2_kb/_0379_ ), .B1(fanout_net_1 ), .B2(\u0_ps2_kb/_0380_ ), .ZN(\u0_ps2_kb/_0381_ ) );
AOI21_X1 \u0_ps2_kb/_0695_ ( .A(\u0_ps2_kb/_0377_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0381_ ), .ZN(\u0_ps2_kb/_0211_ ) );
NOR2_X1 \u0_ps2_kb/_0696_ ( .A1(\u0_ps2_kb/_0347_ ), .A2(\u0_ps2_kb/_0228_ ), .ZN(\u0_ps2_kb/_0382_ ) );
AOI211_X4 \u0_ps2_kb/_0697_ ( .A(\u0_ps2_kb/_0477_ ), .B(\u0_ps2_kb/_0382_ ), .C1(\u0_ps2_kb/_0336_ ), .C2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0383_ ) );
MUX2_X1 \u0_ps2_kb/_0698_ ( .A(\u0_ps2_kb/_0236_ ), .B(\u0_ps2_kb/_0244_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0384_ ) );
AOI211_X4 \u0_ps2_kb/_0699_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0383_ ), .C1(\u0_ps2_kb/_0477_ ), .C2(\u0_ps2_kb/_0384_ ), .ZN(\u0_ps2_kb/_0385_ ) );
MUX2_X1 \u0_ps2_kb/_0700_ ( .A(\u0_ps2_kb/_0252_ ), .B(\u0_ps2_kb/_0268_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0386_ ) );
AND2_X1 \u0_ps2_kb/_0701_ ( .A1(\u0_ps2_kb/_0386_ ), .A2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0387_ ) );
MUX2_X1 \u0_ps2_kb/_0702_ ( .A(\u0_ps2_kb/_0260_ ), .B(\u0_ps2_kb/_0276_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0388_ ) );
AOI21_X1 \u0_ps2_kb/_0703_ ( .A(\u0_ps2_kb/_0387_ ), .B1(fanout_net_1 ), .B2(\u0_ps2_kb/_0388_ ), .ZN(\u0_ps2_kb/_0389_ ) );
AOI21_X1 \u0_ps2_kb/_0704_ ( .A(\u0_ps2_kb/_0385_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0389_ ), .ZN(\u0_ps2_kb/_0212_ ) );
NOR2_X1 \u0_ps2_kb/_0705_ ( .A1(fanout_net_1 ), .A2(\u0_ps2_kb/_0237_ ), .ZN(\u0_ps2_kb/_0390_ ) );
AOI211_X4 \u0_ps2_kb/_0706_ ( .A(\u0_ps2_kb/_0339_ ), .B(\u0_ps2_kb/_0390_ ), .C1(\u0_ps2_kb/_0323_ ), .C2(fanout_net_1 ), .ZN(\u0_ps2_kb/_0391_ ) );
MUX2_X1 \u0_ps2_kb/_0707_ ( .A(\u0_ps2_kb/_0221_ ), .B(\u0_ps2_kb/_0229_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0392_ ) );
AOI211_X4 \u0_ps2_kb/_0708_ ( .A(\u0_ps2_kb/_0478_ ), .B(\u0_ps2_kb/_0391_ ), .C1(\u0_ps2_kb/_0340_ ), .C2(\u0_ps2_kb/_0392_ ), .ZN(\u0_ps2_kb/_0393_ ) );
MUX2_X1 \u0_ps2_kb/_0709_ ( .A(\u0_ps2_kb/_0253_ ), .B(\u0_ps2_kb/_0269_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0394_ ) );
AND2_X1 \u0_ps2_kb/_0710_ ( .A1(\u0_ps2_kb/_0394_ ), .A2(\u0_ps2_kb/_0347_ ), .ZN(\u0_ps2_kb/_0395_ ) );
MUX2_X1 \u0_ps2_kb/_0711_ ( .A(\u0_ps2_kb/_0261_ ), .B(\u0_ps2_kb/_0277_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0396_ ) );
AOI21_X1 \u0_ps2_kb/_0712_ ( .A(\u0_ps2_kb/_0395_ ), .B1(fanout_net_1 ), .B2(\u0_ps2_kb/_0396_ ), .ZN(\u0_ps2_kb/_0397_ ) );
AOI21_X1 \u0_ps2_kb/_0713_ ( .A(\u0_ps2_kb/_0393_ ), .B1(\u0_ps2_kb/_0478_ ), .B2(\u0_ps2_kb/_0397_ ), .ZN(\u0_ps2_kb/_0213_ ) );
MUX2_X1 \u0_ps2_kb/_0714_ ( .A(\u0_ps2_kb/_0222_ ), .B(\u0_ps2_kb/_0238_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0398_ ) );
MUX2_X1 \u0_ps2_kb/_0715_ ( .A(\u0_ps2_kb/_0230_ ), .B(\u0_ps2_kb/_0246_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0399_ ) );
MUX2_X1 \u0_ps2_kb/_0716_ ( .A(\u0_ps2_kb/_0398_ ), .B(\u0_ps2_kb/_0399_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0400_ ) );
MUX2_X1 \u0_ps2_kb/_0717_ ( .A(\u0_ps2_kb/_0254_ ), .B(\u0_ps2_kb/_0270_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0401_ ) );
MUX2_X1 \u0_ps2_kb/_0718_ ( .A(\u0_ps2_kb/_0262_ ), .B(\u0_ps2_kb/_0278_ ), .S(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0402_ ) );
MUX2_X1 \u0_ps2_kb/_0719_ ( .A(\u0_ps2_kb/_0401_ ), .B(\u0_ps2_kb/_0402_ ), .S(fanout_net_1 ), .Z(\u0_ps2_kb/_0403_ ) );
MUX2_X1 \u0_ps2_kb/_0720_ ( .A(\u0_ps2_kb/_0400_ ), .B(\u0_ps2_kb/_0403_ ), .S(\u0_ps2_kb/_0478_ ), .Z(\u0_ps2_kb/_0214_ ) );
INV_X1 \u0_ps2_kb/_0721_ ( .A(\u0_ps2_kb/_0184_ ), .ZN(\u0_ps2_kb/_0404_ ) );
NAND3_X1 \u0_ps2_kb/_0722_ ( .A1(\u0_ps2_kb/_0326_ ), .A2(\u0_ps2_kb/_0404_ ), .A3(\u0_ps2_kb/_0482_ ), .ZN(\u0_ps2_kb/_0405_ ) );
NOR2_X4 \u0_ps2_kb/_0723_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0405_ ), .ZN(\u0_ps2_kb/_0406_ ) );
MUX2_X1 \u0_ps2_kb/_0724_ ( .A(\u0_ps2_kb/_0255_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0158_ ) );
MUX2_X1 \u0_ps2_kb/_0725_ ( .A(\u0_ps2_kb/_0256_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0159_ ) );
MUX2_X1 \u0_ps2_kb/_0726_ ( .A(\u0_ps2_kb/_0257_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0160_ ) );
MUX2_X1 \u0_ps2_kb/_0727_ ( .A(\u0_ps2_kb/_0258_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0161_ ) );
MUX2_X1 \u0_ps2_kb/_0728_ ( .A(\u0_ps2_kb/_0259_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0162_ ) );
MUX2_X1 \u0_ps2_kb/_0729_ ( .A(\u0_ps2_kb/_0260_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0163_ ) );
MUX2_X1 \u0_ps2_kb/_0730_ ( .A(\u0_ps2_kb/_0261_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0164_ ) );
MUX2_X1 \u0_ps2_kb/_0731_ ( .A(\u0_ps2_kb/_0262_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0406_ ), .Z(\u0_ps2_kb/_0165_ ) );
NAND3_X1 \u0_ps2_kb/_0732_ ( .A1(\u0_ps2_kb/_0310_ ), .A2(\u0_ps2_kb/_0326_ ), .A3(\u0_ps2_kb/_0404_ ), .ZN(\u0_ps2_kb/_0407_ ) );
NOR2_X4 \u0_ps2_kb/_0733_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0407_ ), .ZN(\u0_ps2_kb/_0408_ ) );
MUX2_X1 \u0_ps2_kb/_0734_ ( .A(\u0_ps2_kb/_0223_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0126_ ) );
MUX2_X1 \u0_ps2_kb/_0735_ ( .A(\u0_ps2_kb/_0224_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0127_ ) );
MUX2_X1 \u0_ps2_kb/_0736_ ( .A(\u0_ps2_kb/_0225_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0128_ ) );
MUX2_X1 \u0_ps2_kb/_0737_ ( .A(\u0_ps2_kb/_0226_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0129_ ) );
MUX2_X1 \u0_ps2_kb/_0738_ ( .A(\u0_ps2_kb/_0227_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0130_ ) );
MUX2_X1 \u0_ps2_kb/_0739_ ( .A(\u0_ps2_kb/_0228_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0131_ ) );
MUX2_X1 \u0_ps2_kb/_0740_ ( .A(\u0_ps2_kb/_0229_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0132_ ) );
MUX2_X1 \u0_ps2_kb/_0741_ ( .A(\u0_ps2_kb/_0230_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0408_ ), .Z(\u0_ps2_kb/_0133_ ) );
NAND3_X1 \u0_ps2_kb/_0742_ ( .A1(\u0_ps2_kb/_0327_ ), .A2(\u0_ps2_kb/_0482_ ), .A3(\u0_ps2_kb/_0481_ ), .ZN(\u0_ps2_kb/_0409_ ) );
NOR2_X4 \u0_ps2_kb/_0743_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0409_ ), .ZN(\u0_ps2_kb/_0410_ ) );
MUX2_X1 \u0_ps2_kb/_0744_ ( .A(\u0_ps2_kb/_0263_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0166_ ) );
MUX2_X1 \u0_ps2_kb/_0745_ ( .A(\u0_ps2_kb/_0264_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0167_ ) );
MUX2_X1 \u0_ps2_kb/_0746_ ( .A(\u0_ps2_kb/_0265_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0168_ ) );
MUX2_X1 \u0_ps2_kb/_0747_ ( .A(\u0_ps2_kb/_0266_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0169_ ) );
MUX2_X1 \u0_ps2_kb/_0748_ ( .A(\u0_ps2_kb/_0267_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0170_ ) );
MUX2_X1 \u0_ps2_kb/_0749_ ( .A(\u0_ps2_kb/_0268_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0171_ ) );
MUX2_X1 \u0_ps2_kb/_0750_ ( .A(\u0_ps2_kb/_0269_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0172_ ) );
MUX2_X1 \u0_ps2_kb/_0751_ ( .A(\u0_ps2_kb/_0270_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0410_ ), .Z(\u0_ps2_kb/_0173_ ) );
NAND3_X1 \u0_ps2_kb/_0752_ ( .A1(\u0_ps2_kb/_0404_ ), .A2(\u0_ps2_kb/_0482_ ), .A3(\u0_ps2_kb/_0481_ ), .ZN(\u0_ps2_kb/_0411_ ) );
NOR2_X4 \u0_ps2_kb/_0753_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0411_ ), .ZN(\u0_ps2_kb/_0412_ ) );
MUX2_X1 \u0_ps2_kb/_0754_ ( .A(\u0_ps2_kb/_0271_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0174_ ) );
MUX2_X1 \u0_ps2_kb/_0755_ ( .A(\u0_ps2_kb/_0272_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0175_ ) );
MUX2_X1 \u0_ps2_kb/_0756_ ( .A(\u0_ps2_kb/_0273_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0176_ ) );
MUX2_X1 \u0_ps2_kb/_0757_ ( .A(\u0_ps2_kb/_0274_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0177_ ) );
MUX2_X1 \u0_ps2_kb/_0758_ ( .A(\u0_ps2_kb/_0275_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0178_ ) );
MUX2_X1 \u0_ps2_kb/_0759_ ( .A(\u0_ps2_kb/_0276_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0179_ ) );
MUX2_X1 \u0_ps2_kb/_0760_ ( .A(\u0_ps2_kb/_0277_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0180_ ) );
MUX2_X1 \u0_ps2_kb/_0761_ ( .A(\u0_ps2_kb/_0278_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0412_ ), .Z(\u0_ps2_kb/_0181_ ) );
NAND3_X1 \u0_ps2_kb/_0762_ ( .A1(\u0_ps2_kb/_0310_ ), .A2(\u0_ps2_kb/_0327_ ), .A3(\u0_ps2_kb/_0481_ ), .ZN(\u0_ps2_kb/_0413_ ) );
NOR2_X4 \u0_ps2_kb/_0763_ ( .A1(\u0_ps2_kb/_0308_ ), .A2(\u0_ps2_kb/_0413_ ), .ZN(\u0_ps2_kb/_0414_ ) );
MUX2_X1 \u0_ps2_kb/_0764_ ( .A(\u0_ps2_kb/_0231_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0134_ ) );
MUX2_X1 \u0_ps2_kb/_0765_ ( .A(\u0_ps2_kb/_0232_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0135_ ) );
MUX2_X1 \u0_ps2_kb/_0766_ ( .A(\u0_ps2_kb/_0233_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0136_ ) );
MUX2_X1 \u0_ps2_kb/_0767_ ( .A(\u0_ps2_kb/_0234_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0137_ ) );
MUX2_X1 \u0_ps2_kb/_0768_ ( .A(\u0_ps2_kb/_0235_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0138_ ) );
MUX2_X1 \u0_ps2_kb/_0769_ ( .A(\u0_ps2_kb/_0236_ ), .B(\u0_ps2_kb/_0198_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0139_ ) );
MUX2_X1 \u0_ps2_kb/_0770_ ( .A(\u0_ps2_kb/_0237_ ), .B(\u0_ps2_kb/_0199_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0140_ ) );
MUX2_X1 \u0_ps2_kb/_0771_ ( .A(\u0_ps2_kb/_0238_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0414_ ), .Z(\u0_ps2_kb/_0141_ ) );
INV_X1 \u0_ps2_kb/_0772_ ( .A(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0415_ ) );
NOR2_X1 \u0_ps2_kb/_0773_ ( .A1(\u0_ps2_kb/_0415_ ), .A2(\u0_ps2_kb/_0204_ ), .ZN(\u0_ps2_kb/_0416_ ) );
AND2_X1 \u0_ps2_kb/_0774_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0416_ ), .ZN(\u0_ps2_kb/_0417_ ) );
NAND2_X1 \u0_ps2_kb/_0775_ ( .A1(\u0_ps2_kb/_0417_ ), .A2(\u0_ps2_kb/_0287_ ), .ZN(\u0_ps2_kb/_0418_ ) );
MUX2_X1 \u0_ps2_kb/_0776_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0197_ ), .S(\u0_ps2_kb/_0418_ ), .Z(\u0_ps2_kb/_0101_ ) );
AND3_X1 \u0_ps2_kb/_0777_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0415_ ), .A3(\u0_ps2_kb/_0281_ ), .ZN(\u0_ps2_kb/_0419_ ) );
NAND2_X1 \u0_ps2_kb/_0778_ ( .A1(\u0_ps2_kb/_0419_ ), .A2(\u0_ps2_kb/_0287_ ), .ZN(\u0_ps2_kb/_0420_ ) );
MUX2_X1 \u0_ps2_kb/_0779_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0196_ ), .S(\u0_ps2_kb/_0420_ ), .Z(\u0_ps2_kb/_0100_ ) );
NAND2_X1 \u0_ps2_kb/_0780_ ( .A1(\u0_ps2_kb/_0284_ ), .A2(\u0_ps2_kb/_0202_ ), .ZN(\u0_ps2_kb/_0421_ ) );
NOR2_X1 \u0_ps2_kb/_0781_ ( .A1(\u0_ps2_kb/_0421_ ), .A2(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0422_ ) );
NAND2_X1 \u0_ps2_kb/_0782_ ( .A1(\u0_ps2_kb/_0290_ ), .A2(\u0_ps2_kb/_0422_ ), .ZN(\u0_ps2_kb/_0423_ ) );
MUX2_X1 \u0_ps2_kb/_0783_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0195_ ), .S(\u0_ps2_kb/_0423_ ), .Z(\u0_ps2_kb/_0099_ ) );
NAND2_X1 \u0_ps2_kb/_0784_ ( .A1(\u0_ps2_kb/_0283_ ), .A2(\u0_ps2_kb/_0422_ ), .ZN(\u0_ps2_kb/_0424_ ) );
MUX2_X1 \u0_ps2_kb/_0785_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0194_ ), .S(\u0_ps2_kb/_0424_ ), .Z(\u0_ps2_kb/_0098_ ) );
NAND2_X1 \u0_ps2_kb/_0786_ ( .A1(\u0_ps2_kb/_0417_ ), .A2(\u0_ps2_kb/_0422_ ), .ZN(\u0_ps2_kb/_0425_ ) );
MUX2_X1 \u0_ps2_kb/_0787_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0193_ ), .S(\u0_ps2_kb/_0425_ ), .Z(\u0_ps2_kb/_0097_ ) );
NAND2_X1 \u0_ps2_kb/_0788_ ( .A1(\u0_ps2_kb/_0419_ ), .A2(\u0_ps2_kb/_0422_ ), .ZN(\u0_ps2_kb/_0426_ ) );
MUX2_X1 \u0_ps2_kb/_0789_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0192_ ), .S(\u0_ps2_kb/_0426_ ), .Z(\u0_ps2_kb/_0096_ ) );
BUF_X4 \u0_ps2_kb/_0790_ ( .A(\u0_ps2_kb/_0286_ ), .Z(\u0_ps2_kb/_0427_ ) );
XNOR2_X1 \u0_ps2_kb/_0791_ ( .A(\u0_ps2_kb/_0280_ ), .B(\u0_ps2_kb/_0203_ ), .ZN(\u0_ps2_kb/_0428_ ) );
NOR3_X1 \u0_ps2_kb/_0792_ ( .A1(\u0_ps2_kb/_0305_ ), .A2(\u0_ps2_kb/_0427_ ), .A3(\u0_ps2_kb/_0428_ ), .ZN(\u0_ps2_kb/_0106_ ) );
NOR3_X1 \u0_ps2_kb/_0793_ ( .A1(\u0_ps2_kb/_0303_ ), .A2(\u0_ps2_kb/_0203_ ), .A3(\u0_ps2_kb/_0281_ ), .ZN(\u0_ps2_kb/_0429_ ) );
INV_X1 \u0_ps2_kb/_0794_ ( .A(\u0_ps2_kb/_0280_ ), .ZN(\u0_ps2_kb/_0430_ ) );
NOR3_X1 \u0_ps2_kb/_0795_ ( .A1(\u0_ps2_kb/_0429_ ), .A2(\u0_ps2_kb/_0430_ ), .A3(\u0_ps2_kb/_0416_ ), .ZN(\u0_ps2_kb/_0431_ ) );
AOI211_X4 \u0_ps2_kb/_0796_ ( .A(\u0_ps2_kb/_0427_ ), .B(\u0_ps2_kb/_0431_ ), .C1(\u0_ps2_kb/_0185_ ), .C2(\u0_ps2_kb/_0430_ ), .ZN(\u0_ps2_kb/_0107_ ) );
XNOR2_X1 \u0_ps2_kb/_0797_ ( .A(\u0_ps2_kb/_0290_ ), .B(\u0_ps2_kb/_0186_ ), .ZN(\u0_ps2_kb/_0432_ ) );
INV_X1 \u0_ps2_kb/_0798_ ( .A(\u0_ps2_kb/_0305_ ), .ZN(\u0_ps2_kb/_0433_ ) );
AND3_X1 \u0_ps2_kb/_0799_ ( .A1(\u0_ps2_kb/_0432_ ), .A2(\u0_ps2_kb/_0202_ ), .A3(\u0_ps2_kb/_0433_ ), .ZN(\u0_ps2_kb/_0108_ ) );
NAND3_X1 \u0_ps2_kb/_0800_ ( .A1(\u0_ps2_kb/_0280_ ), .A2(\u0_ps2_kb/_0205_ ), .A3(\u0_ps2_kb/_0289_ ), .ZN(\u0_ps2_kb/_0434_ ) );
AOI221_X4 \u0_ps2_kb/_0801_ ( .A(\u0_ps2_kb/_0427_ ), .B1(\u0_ps2_kb/_0434_ ), .B2(\u0_ps2_kb/_0187_ ), .C1(\u0_ps2_kb/_0280_ ), .C2(\u0_ps2_kb/_0304_ ), .ZN(\u0_ps2_kb/_0435_ ) );
OR2_X1 \u0_ps2_kb/_0802_ ( .A1(\u0_ps2_kb/_0434_ ), .A2(\u0_ps2_kb/_0187_ ), .ZN(\u0_ps2_kb/_0436_ ) );
AND2_X1 \u0_ps2_kb/_0803_ ( .A1(\u0_ps2_kb/_0435_ ), .A2(\u0_ps2_kb/_0436_ ), .ZN(\u0_ps2_kb/_0109_ ) );
XOR2_X1 \u0_ps2_kb/_0804_ ( .A(fanout_net_1 ), .B(\u0_ps2_kb/_0471_ ), .Z(\u0_ps2_kb/_0437_ ) );
MUX2_X1 \u0_ps2_kb/_0805_ ( .A(\u0_ps2_kb/_0188_ ), .B(\u0_ps2_kb/_0437_ ), .S(\u0_ps2_kb/_0479_ ), .Z(\u0_ps2_kb/_0438_ ) );
NOR2_X1 \u0_ps2_kb/_0806_ ( .A1(\u0_ps2_kb/_0438_ ), .A2(\u0_ps2_kb/_0427_ ), .ZN(\u0_ps2_kb/_0111_ ) );
XOR2_X1 \u0_ps2_kb/_0807_ ( .A(fanout_net_1 ), .B(\u0_ps2_kb/_0477_ ), .Z(\u0_ps2_kb/_0439_ ) );
INV_X1 \u0_ps2_kb/_0808_ ( .A(\u0_ps2_kb/_0471_ ), .ZN(\u0_ps2_kb/_0440_ ) );
NAND2_X1 \u0_ps2_kb/_0809_ ( .A1(\u0_ps2_kb/_0440_ ), .A2(\u0_ps2_kb/_0479_ ), .ZN(\u0_ps2_kb/_0441_ ) );
NOR2_X1 \u0_ps2_kb/_0810_ ( .A1(\u0_ps2_kb/_0439_ ), .A2(\u0_ps2_kb/_0441_ ), .ZN(\u0_ps2_kb/_0442_ ) );
AOI211_X4 \u0_ps2_kb/_0811_ ( .A(\u0_ps2_kb/_0427_ ), .B(\u0_ps2_kb/_0442_ ), .C1(\u0_ps2_kb/_0183_ ), .C2(\u0_ps2_kb/_0441_ ), .ZN(\u0_ps2_kb/_0112_ ) );
NAND2_X1 \u0_ps2_kb/_0812_ ( .A1(\u0_ps2_kb/_0476_ ), .A2(\u0_ps2_kb/_0477_ ), .ZN(\u0_ps2_kb/_0443_ ) );
XNOR2_X1 \u0_ps2_kb/_0813_ ( .A(\u0_ps2_kb/_0443_ ), .B(\u0_ps2_kb/_0182_ ), .ZN(\u0_ps2_kb/_0444_ ) );
AND3_X1 \u0_ps2_kb/_0814_ ( .A1(\u0_ps2_kb/_0444_ ), .A2(\u0_ps2_kb/_0440_ ), .A3(\u0_ps2_kb/_0479_ ), .ZN(\u0_ps2_kb/_0445_ ) );
AOI211_X4 \u0_ps2_kb/_0815_ ( .A(\u0_ps2_kb/_0427_ ), .B(\u0_ps2_kb/_0445_ ), .C1(\u0_ps2_kb/_0182_ ), .C2(\u0_ps2_kb/_0441_ ), .ZN(\u0_ps2_kb/_0113_ ) );
OAI21_X1 \u0_ps2_kb/_0816_ ( .A(\u0_ps2_kb/_0202_ ), .B1(\u0_ps2_kb/_0306_ ), .B2(\u0_ps2_kb/_0404_ ), .ZN(\u0_ps2_kb/_0446_ ) );
AOI21_X1 \u0_ps2_kb/_0817_ ( .A(\u0_ps2_kb/_0446_ ), .B1(\u0_ps2_kb/_0404_ ), .B2(\u0_ps2_kb/_0306_ ), .ZN(\u0_ps2_kb/_0115_ ) );
AND2_X1 \u0_ps2_kb/_0818_ ( .A1(\u0_ps2_kb/_0302_ ), .A2(\u0_ps2_kb/_0304_ ), .ZN(\u0_ps2_kb/_0447_ ) );
INV_X1 \u0_ps2_kb/_0819_ ( .A(\u0_ps2_kb/_0447_ ), .ZN(\u0_ps2_kb/_0448_ ) );
XNOR2_X1 \u0_ps2_kb/_0820_ ( .A(\u0_ps2_kb/_0481_ ), .B(\u0_ps2_kb/_0480_ ), .ZN(\u0_ps2_kb/_0449_ ) );
NOR2_X2 \u0_ps2_kb/_0821_ ( .A1(\u0_ps2_kb/_0448_ ), .A2(\u0_ps2_kb/_0449_ ), .ZN(\u0_ps2_kb/_0450_ ) );
OAI21_X1 \u0_ps2_kb/_0822_ ( .A(\u0_ps2_kb/_0280_ ), .B1(\u0_ps2_kb/_0447_ ), .B2(\u0_ps2_kb/_0189_ ), .ZN(\u0_ps2_kb/_0451_ ) );
NOR2_X1 \u0_ps2_kb/_0823_ ( .A1(\u0_ps2_kb/_0450_ ), .A2(\u0_ps2_kb/_0451_ ), .ZN(\u0_ps2_kb/_0452_ ) );
AOI211_X2 \u0_ps2_kb/_0824_ ( .A(\u0_ps2_kb/_0427_ ), .B(\u0_ps2_kb/_0452_ ), .C1(\u0_ps2_kb/_0189_ ), .C2(\u0_ps2_kb/_0430_ ), .ZN(\u0_ps2_kb/_0116_ ) );
NAND2_X1 \u0_ps2_kb/_0825_ ( .A1(\u0_ps2_kb/_0481_ ), .A2(\u0_ps2_kb/_0480_ ), .ZN(\u0_ps2_kb/_0453_ ) );
XNOR2_X1 \u0_ps2_kb/_0826_ ( .A(\u0_ps2_kb/_0453_ ), .B(\u0_ps2_kb/_0190_ ), .ZN(\u0_ps2_kb/_0454_ ) );
AND4_X1 \u0_ps2_kb/_0827_ ( .A1(\u0_ps2_kb/_0301_ ), .A2(\u0_ps2_kb/_0300_ ), .A3(\u0_ps2_kb/_0305_ ), .A4(\u0_ps2_kb/_0454_ ), .ZN(\u0_ps2_kb/_0455_ ) );
INV_X1 \u0_ps2_kb/_0828_ ( .A(\u0_ps2_kb/_0306_ ), .ZN(\u0_ps2_kb/_0456_ ) );
AOI211_X4 \u0_ps2_kb/_0829_ ( .A(\u0_ps2_kb/_0427_ ), .B(\u0_ps2_kb/_0455_ ), .C1(\u0_ps2_kb/_0456_ ), .C2(\u0_ps2_kb/_0190_ ), .ZN(\u0_ps2_kb/_0117_ ) );
NOR3_X1 \u0_ps2_kb/_0830_ ( .A1(\u0_ps2_kb/_0427_ ), .A2(\u0_ps2_kb/_0284_ ), .A3(\u0_ps2_kb/_0205_ ), .ZN(\u0_ps2_kb/_0457_ ) );
NAND2_X1 \u0_ps2_kb/_0831_ ( .A1(\u0_ps2_kb/_0419_ ), .A2(\u0_ps2_kb/_0457_ ), .ZN(\u0_ps2_kb/_0458_ ) );
MUX2_X1 \u0_ps2_kb/_0832_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0200_ ), .S(\u0_ps2_kb/_0458_ ), .Z(\u0_ps2_kb/_0104_ ) );
NAND2_X1 \u0_ps2_kb/_0833_ ( .A1(\u0_ps2_kb/_0417_ ), .A2(\u0_ps2_kb/_0457_ ), .ZN(\u0_ps2_kb/_0459_ ) );
MUX2_X1 \u0_ps2_kb/_0834_ ( .A(\u0_ps2_kb/_0475_ ), .B(\u0_ps2_kb/_0201_ ), .S(\u0_ps2_kb/_0459_ ), .Z(\u0_ps2_kb/_0105_ ) );
XOR2_X1 \u0_ps2_kb/_0835_ ( .A(\u0_ps2_kb/_0439_ ), .B(\u0_ps2_kb/_0189_ ), .Z(\u0_ps2_kb/_0460_ ) );
XNOR2_X1 \u0_ps2_kb/_0836_ ( .A(\u0_ps2_kb/_0444_ ), .B(\u0_ps2_kb/_0190_ ), .ZN(\u0_ps2_kb/_0461_ ) );
XNOR2_X1 \u0_ps2_kb/_0837_ ( .A(\u0_ps2_kb/_0480_ ), .B(\u0_ps2_kb/_0476_ ), .ZN(\u0_ps2_kb/_0462_ ) );
NOR2_X1 \u0_ps2_kb/_0838_ ( .A1(\u0_ps2_kb/_0462_ ), .A2(\u0_ps2_kb/_0471_ ), .ZN(\u0_ps2_kb/_0463_ ) );
NAND3_X1 \u0_ps2_kb/_0839_ ( .A1(\u0_ps2_kb/_0460_ ), .A2(\u0_ps2_kb/_0461_ ), .A3(\u0_ps2_kb/_0463_ ), .ZN(\u0_ps2_kb/_0464_ ) );
NAND3_X1 \u0_ps2_kb/_0840_ ( .A1(\u0_ps2_kb/_0464_ ), .A2(\u0_ps2_kb/_0202_ ), .A3(\u0_ps2_kb/_0479_ ), .ZN(\u0_ps2_kb/_0465_ ) );
NAND2_X1 \u0_ps2_kb/_0841_ ( .A1(\u0_ps2_kb/_0309_ ), .A2(\u0_ps2_kb/_0465_ ), .ZN(\u0_ps2_kb/_0114_ ) );
XOR2_X1 \u0_ps2_kb/_0842_ ( .A(\u0_ps2_kb/_0454_ ), .B(\u0_ps2_kb/_0182_ ), .Z(\u0_ps2_kb/_0466_ ) );
XOR2_X1 \u0_ps2_kb/_0843_ ( .A(\u0_ps2_kb/_0449_ ), .B(\u0_ps2_kb/_0183_ ), .Z(\u0_ps2_kb/_0467_ ) );
NOR3_X1 \u0_ps2_kb/_0844_ ( .A1(\u0_ps2_kb/_0466_ ), .A2(\u0_ps2_kb/_0462_ ), .A3(\u0_ps2_kb/_0467_ ), .ZN(\u0_ps2_kb/_0468_ ) );
NAND3_X1 \u0_ps2_kb/_0845_ ( .A1(\u0_ps2_kb/_0300_ ), .A2(\u0_ps2_kb/_0301_ ), .A3(\u0_ps2_kb/_0468_ ), .ZN(\u0_ps2_kb/_0469_ ) );
NOR2_X1 \u0_ps2_kb/_0846_ ( .A1(\u0_ps2_kb/_0433_ ), .A2(\u0_ps2_kb/_0472_ ), .ZN(\u0_ps2_kb/_0470_ ) );
AOI221_X4 \u0_ps2_kb/_0847_ ( .A(\u0_ps2_kb/_0427_ ), .B1(\u0_ps2_kb/_0191_ ), .B2(\u0_ps2_kb/_0433_ ), .C1(\u0_ps2_kb/_0469_ ), .C2(\u0_ps2_kb/_0470_ ), .ZN(\u0_ps2_kb/_0110_ ) );
BUF_X1 \u0_ps2_kb/_0848_ ( .A(fanout_net_2 ), .Z(\u0_ps2_kb/_0202_ ) );
BUF_X1 \u0_ps2_kb/_0849_ ( .A(\u0_ps2_kb/ps2_clk_sync[1] ), .Z(\u0_ps2_kb/_0473_ ) );
BUF_X1 \u0_ps2_kb/_0850_ ( .A(\u0_ps2_kb/ps2_clk_sync[2] ), .Z(\u0_ps2_kb/_0474_ ) );
BUF_X1 \u0_ps2_kb/_0851_ ( .A(\u0_ps2_kb/count[0] ), .Z(\u0_ps2_kb/_0203_ ) );
BUF_X1 \u0_ps2_kb/_0852_ ( .A(\u0_ps2_kb/count[1] ), .Z(\u0_ps2_kb/_0204_ ) );
BUF_X1 \u0_ps2_kb/_0853_ ( .A(\u0_ps2_kb/count[2] ), .Z(\u0_ps2_kb/_0205_ ) );
BUF_X1 \u0_ps2_kb/_0854_ ( .A(\u0_ps2_kb/count[3] ), .Z(\u0_ps2_kb/_0206_ ) );
BUF_X1 \u0_ps2_kb/_0855_ ( .A(ps2_data ), .Z(\u0_ps2_kb/_0475_ ) );
BUF_X1 \u0_ps2_kb/_0856_ ( .A(\u0_ps2_kb/buffer[6] ), .Z(\u0_ps2_kb/_0198_ ) );
BUF_X1 \u0_ps2_kb/_0857_ ( .A(\u0_ps2_kb/_0102_ ), .Z(\u0_ps2_kb/_0006_ ) );
BUF_X1 \u0_ps2_kb/_0858_ ( .A(\u0_ps2_kb/buffer[7] ), .Z(\u0_ps2_kb/_0199_ ) );
BUF_X1 \u0_ps2_kb/_0859_ ( .A(\u0_ps2_kb/_0103_ ), .Z(\u0_ps2_kb/_0007_ ) );
BUF_X1 \u0_ps2_kb/_0860_ ( .A(\u0_ps2_kb/w_ptr[2] ), .Z(\u0_ps2_kb/_0482_ ) );
BUF_X1 \u0_ps2_kb/_0861_ ( .A(\u0_ps2_kb/w_ptr[1] ), .Z(\u0_ps2_kb/_0481_ ) );
BUF_X1 \u0_ps2_kb/_0862_ ( .A(\u0_ps2_kb/w_ptr[0] ), .Z(\u0_ps2_kb/_0480_ ) );
BUF_X1 \u0_ps2_kb/_0863_ ( .A(\u0_ps2_kb/buffer[0] ), .Z(\u0_ps2_kb/_0192_ ) );
BUF_X1 \u0_ps2_kb/_0864_ ( .A(\u0_ps2_kb/buffer[2] ), .Z(\u0_ps2_kb/_0194_ ) );
BUF_X1 \u0_ps2_kb/_0865_ ( .A(\u0_ps2_kb/buffer[1] ), .Z(\u0_ps2_kb/_0193_ ) );
BUF_X1 \u0_ps2_kb/_0866_ ( .A(\u0_ps2_kb/buffer[4] ), .Z(\u0_ps2_kb/_0196_ ) );
BUF_X1 \u0_ps2_kb/_0867_ ( .A(\u0_ps2_kb/buffer[3] ), .Z(\u0_ps2_kb/_0195_ ) );
BUF_X1 \u0_ps2_kb/_0868_ ( .A(\u0_ps2_kb/buffer[5] ), .Z(\u0_ps2_kb/_0197_ ) );
BUF_X1 \u0_ps2_kb/_0869_ ( .A(\u0_ps2_kb/buffer[8] ), .Z(\u0_ps2_kb/_0200_ ) );
BUF_X1 \u0_ps2_kb/_0870_ ( .A(\u0_ps2_kb/buffer[9] ), .Z(\u0_ps2_kb/_0201_ ) );
BUF_X1 \u0_ps2_kb/_0871_ ( .A(\u0_ps2_kb/fifo[3][0] ), .Z(\u0_ps2_kb/_0239_ ) );
BUF_X1 \u0_ps2_kb/_0872_ ( .A(\u0_ps2_kb/_0142_ ), .Z(\u0_ps2_kb/_0046_ ) );
BUF_X1 \u0_ps2_kb/_0873_ ( .A(\u0_ps2_kb/fifo[3][1] ), .Z(\u0_ps2_kb/_0240_ ) );
BUF_X1 \u0_ps2_kb/_0874_ ( .A(\u0_ps2_kb/_0143_ ), .Z(\u0_ps2_kb/_0047_ ) );
BUF_X1 \u0_ps2_kb/_0875_ ( .A(\u0_ps2_kb/fifo[3][2] ), .Z(\u0_ps2_kb/_0241_ ) );
BUF_X1 \u0_ps2_kb/_0876_ ( .A(\u0_ps2_kb/_0144_ ), .Z(\u0_ps2_kb/_0048_ ) );
BUF_X1 \u0_ps2_kb/_0877_ ( .A(\u0_ps2_kb/fifo[3][3] ), .Z(\u0_ps2_kb/_0242_ ) );
BUF_X1 \u0_ps2_kb/_0878_ ( .A(\u0_ps2_kb/_0145_ ), .Z(\u0_ps2_kb/_0049_ ) );
BUF_X1 \u0_ps2_kb/_0879_ ( .A(\u0_ps2_kb/fifo[3][4] ), .Z(\u0_ps2_kb/_0243_ ) );
BUF_X1 \u0_ps2_kb/_0880_ ( .A(\u0_ps2_kb/_0146_ ), .Z(\u0_ps2_kb/_0050_ ) );
BUF_X1 \u0_ps2_kb/_0881_ ( .A(\u0_ps2_kb/fifo[3][5] ), .Z(\u0_ps2_kb/_0244_ ) );
BUF_X1 \u0_ps2_kb/_0882_ ( .A(\u0_ps2_kb/_0147_ ), .Z(\u0_ps2_kb/_0051_ ) );
BUF_X1 \u0_ps2_kb/_0883_ ( .A(\u0_ps2_kb/fifo[3][6] ), .Z(\u0_ps2_kb/_0245_ ) );
BUF_X1 \u0_ps2_kb/_0884_ ( .A(\u0_ps2_kb/_0148_ ), .Z(\u0_ps2_kb/_0052_ ) );
BUF_X1 \u0_ps2_kb/_0885_ ( .A(\u0_ps2_kb/fifo[3][7] ), .Z(\u0_ps2_kb/_0246_ ) );
BUF_X1 \u0_ps2_kb/_0886_ ( .A(\u0_ps2_kb/_0149_ ), .Z(\u0_ps2_kb/_0053_ ) );
BUF_X1 \u0_ps2_kb/_0887_ ( .A(\u0_ps2_kb/fifo[4][0] ), .Z(\u0_ps2_kb/_0247_ ) );
BUF_X1 \u0_ps2_kb/_0888_ ( .A(\u0_ps2_kb/_0150_ ), .Z(\u0_ps2_kb/_0054_ ) );
BUF_X1 \u0_ps2_kb/_0889_ ( .A(\u0_ps2_kb/fifo[4][1] ), .Z(\u0_ps2_kb/_0248_ ) );
BUF_X1 \u0_ps2_kb/_0890_ ( .A(\u0_ps2_kb/_0151_ ), .Z(\u0_ps2_kb/_0055_ ) );
BUF_X1 \u0_ps2_kb/_0891_ ( .A(\u0_ps2_kb/fifo[4][2] ), .Z(\u0_ps2_kb/_0249_ ) );
BUF_X1 \u0_ps2_kb/_0892_ ( .A(\u0_ps2_kb/_0152_ ), .Z(\u0_ps2_kb/_0056_ ) );
BUF_X1 \u0_ps2_kb/_0893_ ( .A(\u0_ps2_kb/fifo[4][3] ), .Z(\u0_ps2_kb/_0250_ ) );
BUF_X1 \u0_ps2_kb/_0894_ ( .A(\u0_ps2_kb/_0153_ ), .Z(\u0_ps2_kb/_0057_ ) );
BUF_X1 \u0_ps2_kb/_0895_ ( .A(\u0_ps2_kb/fifo[4][4] ), .Z(\u0_ps2_kb/_0251_ ) );
BUF_X1 \u0_ps2_kb/_0896_ ( .A(\u0_ps2_kb/_0154_ ), .Z(\u0_ps2_kb/_0058_ ) );
BUF_X1 \u0_ps2_kb/_0897_ ( .A(\u0_ps2_kb/fifo[4][5] ), .Z(\u0_ps2_kb/_0252_ ) );
BUF_X1 \u0_ps2_kb/_0898_ ( .A(\u0_ps2_kb/_0155_ ), .Z(\u0_ps2_kb/_0059_ ) );
BUF_X1 \u0_ps2_kb/_0899_ ( .A(\u0_ps2_kb/fifo[4][6] ), .Z(\u0_ps2_kb/_0253_ ) );
BUF_X1 \u0_ps2_kb/_0900_ ( .A(\u0_ps2_kb/_0156_ ), .Z(\u0_ps2_kb/_0060_ ) );
BUF_X1 \u0_ps2_kb/_0901_ ( .A(\u0_ps2_kb/fifo[4][7] ), .Z(\u0_ps2_kb/_0254_ ) );
BUF_X1 \u0_ps2_kb/_0902_ ( .A(\u0_ps2_kb/_0157_ ), .Z(\u0_ps2_kb/_0061_ ) );
BUF_X1 \u0_ps2_kb/_0903_ ( .A(\u0_ps2_kb/fifo[0][0] ), .Z(\u0_ps2_kb/_0215_ ) );
BUF_X1 \u0_ps2_kb/_0904_ ( .A(\u0_ps2_kb/_0118_ ), .Z(\u0_ps2_kb/_0022_ ) );
BUF_X1 \u0_ps2_kb/_0905_ ( .A(\u0_ps2_kb/fifo[0][1] ), .Z(\u0_ps2_kb/_0216_ ) );
BUF_X1 \u0_ps2_kb/_0906_ ( .A(\u0_ps2_kb/_0119_ ), .Z(\u0_ps2_kb/_0023_ ) );
BUF_X1 \u0_ps2_kb/_0907_ ( .A(\u0_ps2_kb/fifo[0][2] ), .Z(\u0_ps2_kb/_0217_ ) );
BUF_X1 \u0_ps2_kb/_0908_ ( .A(\u0_ps2_kb/_0120_ ), .Z(\u0_ps2_kb/_0024_ ) );
BUF_X1 \u0_ps2_kb/_0909_ ( .A(\u0_ps2_kb/fifo[0][3] ), .Z(\u0_ps2_kb/_0218_ ) );
BUF_X1 \u0_ps2_kb/_0910_ ( .A(\u0_ps2_kb/_0121_ ), .Z(\u0_ps2_kb/_0025_ ) );
BUF_X1 \u0_ps2_kb/_0911_ ( .A(\u0_ps2_kb/fifo[0][4] ), .Z(\u0_ps2_kb/_0219_ ) );
BUF_X1 \u0_ps2_kb/_0912_ ( .A(\u0_ps2_kb/_0122_ ), .Z(\u0_ps2_kb/_0026_ ) );
BUF_X1 \u0_ps2_kb/_0913_ ( .A(\u0_ps2_kb/fifo[0][5] ), .Z(\u0_ps2_kb/_0220_ ) );
BUF_X1 \u0_ps2_kb/_0914_ ( .A(\u0_ps2_kb/_0123_ ), .Z(\u0_ps2_kb/_0027_ ) );
BUF_X1 \u0_ps2_kb/_0915_ ( .A(\u0_ps2_kb/fifo[0][6] ), .Z(\u0_ps2_kb/_0221_ ) );
BUF_X1 \u0_ps2_kb/_0916_ ( .A(\u0_ps2_kb/_0124_ ), .Z(\u0_ps2_kb/_0028_ ) );
BUF_X1 \u0_ps2_kb/_0917_ ( .A(\u0_ps2_kb/fifo[0][7] ), .Z(\u0_ps2_kb/_0222_ ) );
BUF_X1 \u0_ps2_kb/_0918_ ( .A(\u0_ps2_kb/_0125_ ), .Z(\u0_ps2_kb/_0029_ ) );
BUF_X1 \u0_ps2_kb/_0919_ ( .A(\u0_ps2_kb/fifo[1][0] ), .Z(\u0_ps2_kb/_0223_ ) );
BUF_X1 \u0_ps2_kb/_0920_ ( .A(\u0_ps2_kb/r_ptr[0] ), .Z(\u0_ps2_kb/_0476_ ) );
BUF_X1 \u0_ps2_kb/_0921_ ( .A(\u0_ps2_kb/fifo[2][0] ), .Z(\u0_ps2_kb/_0231_ ) );
BUF_X1 \u0_ps2_kb/_0922_ ( .A(\u0_ps2_kb/r_ptr[1] ), .Z(\u0_ps2_kb/_0477_ ) );
BUF_X1 \u0_ps2_kb/_0923_ ( .A(\u0_ps2_kb/fifo[5][0] ), .Z(\u0_ps2_kb/_0255_ ) );
BUF_X1 \u0_ps2_kb/_0924_ ( .A(\u0_ps2_kb/fifo[6][0] ), .Z(\u0_ps2_kb/_0263_ ) );
BUF_X1 \u0_ps2_kb/_0925_ ( .A(\u0_ps2_kb/fifo[7][0] ), .Z(\u0_ps2_kb/_0271_ ) );
BUF_X1 \u0_ps2_kb/_0926_ ( .A(\u0_ps2_kb/r_ptr[2] ), .Z(\u0_ps2_kb/_0478_ ) );
BUF_X1 \u0_ps2_kb/_0927_ ( .A(\u0_ps2_kb/_0207_ ), .Z(\data[0] ) );
BUF_X1 \u0_ps2_kb/_0928_ ( .A(\u0_ps2_kb/fifo[1][1] ), .Z(\u0_ps2_kb/_0224_ ) );
BUF_X1 \u0_ps2_kb/_0929_ ( .A(\u0_ps2_kb/fifo[2][1] ), .Z(\u0_ps2_kb/_0232_ ) );
BUF_X1 \u0_ps2_kb/_0930_ ( .A(\u0_ps2_kb/fifo[5][1] ), .Z(\u0_ps2_kb/_0256_ ) );
BUF_X1 \u0_ps2_kb/_0931_ ( .A(\u0_ps2_kb/fifo[6][1] ), .Z(\u0_ps2_kb/_0264_ ) );
BUF_X1 \u0_ps2_kb/_0932_ ( .A(\u0_ps2_kb/fifo[7][1] ), .Z(\u0_ps2_kb/_0272_ ) );
BUF_X1 \u0_ps2_kb/_0933_ ( .A(\u0_ps2_kb/_0208_ ), .Z(\data[1] ) );
BUF_X1 \u0_ps2_kb/_0934_ ( .A(\u0_ps2_kb/fifo[1][2] ), .Z(\u0_ps2_kb/_0225_ ) );
BUF_X1 \u0_ps2_kb/_0935_ ( .A(\u0_ps2_kb/fifo[2][2] ), .Z(\u0_ps2_kb/_0233_ ) );
BUF_X1 \u0_ps2_kb/_0936_ ( .A(\u0_ps2_kb/fifo[5][2] ), .Z(\u0_ps2_kb/_0257_ ) );
BUF_X1 \u0_ps2_kb/_0937_ ( .A(\u0_ps2_kb/fifo[6][2] ), .Z(\u0_ps2_kb/_0265_ ) );
BUF_X1 \u0_ps2_kb/_0938_ ( .A(\u0_ps2_kb/fifo[7][2] ), .Z(\u0_ps2_kb/_0273_ ) );
BUF_X1 \u0_ps2_kb/_0939_ ( .A(\u0_ps2_kb/_0209_ ), .Z(\data[2] ) );
BUF_X1 \u0_ps2_kb/_0940_ ( .A(\u0_ps2_kb/fifo[1][3] ), .Z(\u0_ps2_kb/_0226_ ) );
BUF_X1 \u0_ps2_kb/_0941_ ( .A(\u0_ps2_kb/fifo[2][3] ), .Z(\u0_ps2_kb/_0234_ ) );
BUF_X1 \u0_ps2_kb/_0942_ ( .A(\u0_ps2_kb/fifo[5][3] ), .Z(\u0_ps2_kb/_0258_ ) );
BUF_X1 \u0_ps2_kb/_0943_ ( .A(\u0_ps2_kb/fifo[6][3] ), .Z(\u0_ps2_kb/_0266_ ) );
BUF_X1 \u0_ps2_kb/_0944_ ( .A(\u0_ps2_kb/fifo[7][3] ), .Z(\u0_ps2_kb/_0274_ ) );
BUF_X1 \u0_ps2_kb/_0945_ ( .A(\u0_ps2_kb/_0210_ ), .Z(\data[3] ) );
BUF_X1 \u0_ps2_kb/_0946_ ( .A(\u0_ps2_kb/fifo[1][4] ), .Z(\u0_ps2_kb/_0227_ ) );
BUF_X1 \u0_ps2_kb/_0947_ ( .A(\u0_ps2_kb/fifo[2][4] ), .Z(\u0_ps2_kb/_0235_ ) );
BUF_X1 \u0_ps2_kb/_0948_ ( .A(\u0_ps2_kb/fifo[5][4] ), .Z(\u0_ps2_kb/_0259_ ) );
BUF_X1 \u0_ps2_kb/_0949_ ( .A(\u0_ps2_kb/fifo[6][4] ), .Z(\u0_ps2_kb/_0267_ ) );
BUF_X1 \u0_ps2_kb/_0950_ ( .A(\u0_ps2_kb/fifo[7][4] ), .Z(\u0_ps2_kb/_0275_ ) );
BUF_X1 \u0_ps2_kb/_0951_ ( .A(\u0_ps2_kb/_0211_ ), .Z(\data[4] ) );
BUF_X1 \u0_ps2_kb/_0952_ ( .A(\u0_ps2_kb/fifo[1][5] ), .Z(\u0_ps2_kb/_0228_ ) );
BUF_X1 \u0_ps2_kb/_0953_ ( .A(\u0_ps2_kb/fifo[2][5] ), .Z(\u0_ps2_kb/_0236_ ) );
BUF_X1 \u0_ps2_kb/_0954_ ( .A(\u0_ps2_kb/fifo[5][5] ), .Z(\u0_ps2_kb/_0260_ ) );
BUF_X1 \u0_ps2_kb/_0955_ ( .A(\u0_ps2_kb/fifo[6][5] ), .Z(\u0_ps2_kb/_0268_ ) );
BUF_X1 \u0_ps2_kb/_0956_ ( .A(\u0_ps2_kb/fifo[7][5] ), .Z(\u0_ps2_kb/_0276_ ) );
BUF_X1 \u0_ps2_kb/_0957_ ( .A(\u0_ps2_kb/_0212_ ), .Z(\data[5] ) );
BUF_X1 \u0_ps2_kb/_0958_ ( .A(\u0_ps2_kb/fifo[1][6] ), .Z(\u0_ps2_kb/_0229_ ) );
BUF_X1 \u0_ps2_kb/_0959_ ( .A(\u0_ps2_kb/fifo[2][6] ), .Z(\u0_ps2_kb/_0237_ ) );
BUF_X1 \u0_ps2_kb/_0960_ ( .A(\u0_ps2_kb/fifo[5][6] ), .Z(\u0_ps2_kb/_0261_ ) );
BUF_X1 \u0_ps2_kb/_0961_ ( .A(\u0_ps2_kb/fifo[6][6] ), .Z(\u0_ps2_kb/_0269_ ) );
BUF_X1 \u0_ps2_kb/_0962_ ( .A(\u0_ps2_kb/fifo[7][6] ), .Z(\u0_ps2_kb/_0277_ ) );
BUF_X1 \u0_ps2_kb/_0963_ ( .A(\u0_ps2_kb/_0213_ ), .Z(\data[6] ) );
BUF_X1 \u0_ps2_kb/_0964_ ( .A(\u0_ps2_kb/fifo[1][7] ), .Z(\u0_ps2_kb/_0230_ ) );
BUF_X1 \u0_ps2_kb/_0965_ ( .A(\u0_ps2_kb/fifo[2][7] ), .Z(\u0_ps2_kb/_0238_ ) );
BUF_X1 \u0_ps2_kb/_0966_ ( .A(\u0_ps2_kb/fifo[5][7] ), .Z(\u0_ps2_kb/_0262_ ) );
BUF_X1 \u0_ps2_kb/_0967_ ( .A(\u0_ps2_kb/fifo[6][7] ), .Z(\u0_ps2_kb/_0270_ ) );
BUF_X1 \u0_ps2_kb/_0968_ ( .A(\u0_ps2_kb/fifo[7][7] ), .Z(\u0_ps2_kb/_0278_ ) );
BUF_X1 \u0_ps2_kb/_0969_ ( .A(\u0_ps2_kb/_0214_ ), .Z(\data[7] ) );
BUF_X1 \u0_ps2_kb/_0970_ ( .A(\u0_ps2_kb/_0088_ ), .Z(\u0_ps2_kb/_0184_ ) );
BUF_X1 \u0_ps2_kb/_0971_ ( .A(\u0_ps2_kb/_0158_ ), .Z(\u0_ps2_kb/_0062_ ) );
BUF_X1 \u0_ps2_kb/_0972_ ( .A(\u0_ps2_kb/_0159_ ), .Z(\u0_ps2_kb/_0063_ ) );
BUF_X1 \u0_ps2_kb/_0973_ ( .A(\u0_ps2_kb/_0160_ ), .Z(\u0_ps2_kb/_0064_ ) );
BUF_X1 \u0_ps2_kb/_0974_ ( .A(\u0_ps2_kb/_0161_ ), .Z(\u0_ps2_kb/_0065_ ) );
BUF_X1 \u0_ps2_kb/_0975_ ( .A(\u0_ps2_kb/_0162_ ), .Z(\u0_ps2_kb/_0066_ ) );
BUF_X1 \u0_ps2_kb/_0976_ ( .A(\u0_ps2_kb/_0163_ ), .Z(\u0_ps2_kb/_0067_ ) );
BUF_X1 \u0_ps2_kb/_0977_ ( .A(\u0_ps2_kb/_0164_ ), .Z(\u0_ps2_kb/_0068_ ) );
BUF_X1 \u0_ps2_kb/_0978_ ( .A(\u0_ps2_kb/_0165_ ), .Z(\u0_ps2_kb/_0069_ ) );
BUF_X1 \u0_ps2_kb/_0979_ ( .A(\u0_ps2_kb/_0126_ ), .Z(\u0_ps2_kb/_0030_ ) );
BUF_X1 \u0_ps2_kb/_0980_ ( .A(\u0_ps2_kb/_0127_ ), .Z(\u0_ps2_kb/_0031_ ) );
BUF_X1 \u0_ps2_kb/_0981_ ( .A(\u0_ps2_kb/_0128_ ), .Z(\u0_ps2_kb/_0032_ ) );
BUF_X1 \u0_ps2_kb/_0982_ ( .A(\u0_ps2_kb/_0129_ ), .Z(\u0_ps2_kb/_0033_ ) );
BUF_X1 \u0_ps2_kb/_0983_ ( .A(\u0_ps2_kb/_0130_ ), .Z(\u0_ps2_kb/_0034_ ) );
BUF_X1 \u0_ps2_kb/_0984_ ( .A(\u0_ps2_kb/_0131_ ), .Z(\u0_ps2_kb/_0035_ ) );
BUF_X1 \u0_ps2_kb/_0985_ ( .A(\u0_ps2_kb/_0132_ ), .Z(\u0_ps2_kb/_0036_ ) );
BUF_X1 \u0_ps2_kb/_0986_ ( .A(\u0_ps2_kb/_0133_ ), .Z(\u0_ps2_kb/_0037_ ) );
BUF_X1 \u0_ps2_kb/_0987_ ( .A(\u0_ps2_kb/_0166_ ), .Z(\u0_ps2_kb/_0070_ ) );
BUF_X1 \u0_ps2_kb/_0988_ ( .A(\u0_ps2_kb/_0167_ ), .Z(\u0_ps2_kb/_0071_ ) );
BUF_X1 \u0_ps2_kb/_0989_ ( .A(\u0_ps2_kb/_0168_ ), .Z(\u0_ps2_kb/_0072_ ) );
BUF_X1 \u0_ps2_kb/_0990_ ( .A(\u0_ps2_kb/_0169_ ), .Z(\u0_ps2_kb/_0073_ ) );
BUF_X1 \u0_ps2_kb/_0991_ ( .A(\u0_ps2_kb/_0170_ ), .Z(\u0_ps2_kb/_0074_ ) );
BUF_X1 \u0_ps2_kb/_0992_ ( .A(\u0_ps2_kb/_0171_ ), .Z(\u0_ps2_kb/_0075_ ) );
BUF_X1 \u0_ps2_kb/_0993_ ( .A(\u0_ps2_kb/_0172_ ), .Z(\u0_ps2_kb/_0076_ ) );
BUF_X1 \u0_ps2_kb/_0994_ ( .A(\u0_ps2_kb/_0173_ ), .Z(\u0_ps2_kb/_0077_ ) );
BUF_X1 \u0_ps2_kb/_0995_ ( .A(\u0_ps2_kb/_0174_ ), .Z(\u0_ps2_kb/_0078_ ) );
BUF_X1 \u0_ps2_kb/_0996_ ( .A(\u0_ps2_kb/_0175_ ), .Z(\u0_ps2_kb/_0079_ ) );
BUF_X1 \u0_ps2_kb/_0997_ ( .A(\u0_ps2_kb/_0176_ ), .Z(\u0_ps2_kb/_0080_ ) );
BUF_X1 \u0_ps2_kb/_0998_ ( .A(\u0_ps2_kb/_0177_ ), .Z(\u0_ps2_kb/_0081_ ) );
BUF_X1 \u0_ps2_kb/_0999_ ( .A(\u0_ps2_kb/_0178_ ), .Z(\u0_ps2_kb/_0082_ ) );
BUF_X1 \u0_ps2_kb/_1000_ ( .A(\u0_ps2_kb/_0179_ ), .Z(\u0_ps2_kb/_0083_ ) );
BUF_X1 \u0_ps2_kb/_1001_ ( .A(\u0_ps2_kb/_0180_ ), .Z(\u0_ps2_kb/_0084_ ) );
BUF_X1 \u0_ps2_kb/_1002_ ( .A(\u0_ps2_kb/_0181_ ), .Z(\u0_ps2_kb/_0085_ ) );
BUF_X1 \u0_ps2_kb/_1003_ ( .A(\u0_ps2_kb/_0134_ ), .Z(\u0_ps2_kb/_0038_ ) );
BUF_X1 \u0_ps2_kb/_1004_ ( .A(\u0_ps2_kb/_0135_ ), .Z(\u0_ps2_kb/_0039_ ) );
BUF_X1 \u0_ps2_kb/_1005_ ( .A(\u0_ps2_kb/_0136_ ), .Z(\u0_ps2_kb/_0040_ ) );
BUF_X1 \u0_ps2_kb/_1006_ ( .A(\u0_ps2_kb/_0137_ ), .Z(\u0_ps2_kb/_0041_ ) );
BUF_X1 \u0_ps2_kb/_1007_ ( .A(\u0_ps2_kb/_0138_ ), .Z(\u0_ps2_kb/_0042_ ) );
BUF_X1 \u0_ps2_kb/_1008_ ( .A(\u0_ps2_kb/_0139_ ), .Z(\u0_ps2_kb/_0043_ ) );
BUF_X1 \u0_ps2_kb/_1009_ ( .A(\u0_ps2_kb/_0140_ ), .Z(\u0_ps2_kb/_0044_ ) );
BUF_X1 \u0_ps2_kb/_1010_ ( .A(\u0_ps2_kb/_0141_ ), .Z(\u0_ps2_kb/_0045_ ) );
BUF_X1 \u0_ps2_kb/_1011_ ( .A(\u0_ps2_kb/_0101_ ), .Z(\u0_ps2_kb/_0005_ ) );
BUF_X1 \u0_ps2_kb/_1012_ ( .A(\u0_ps2_kb/_0100_ ), .Z(\u0_ps2_kb/_0004_ ) );
BUF_X1 \u0_ps2_kb/_1013_ ( .A(\u0_ps2_kb/_0099_ ), .Z(\u0_ps2_kb/_0003_ ) );
BUF_X1 \u0_ps2_kb/_1014_ ( .A(\u0_ps2_kb/_0098_ ), .Z(\u0_ps2_kb/_0002_ ) );
BUF_X1 \u0_ps2_kb/_1015_ ( .A(\u0_ps2_kb/_0097_ ), .Z(\u0_ps2_kb/_0001_ ) );
BUF_X1 \u0_ps2_kb/_1016_ ( .A(\u0_ps2_kb/_0096_ ), .Z(\u0_ps2_kb/_0000_ ) );
BUF_X1 \u0_ps2_kb/_1017_ ( .A(\u0_ps2_kb/_0106_ ), .Z(\u0_ps2_kb/_0010_ ) );
BUF_X1 \u0_ps2_kb/_1018_ ( .A(\u0_ps2_kb/_0089_ ), .Z(\u0_ps2_kb/_0185_ ) );
BUF_X1 \u0_ps2_kb/_1019_ ( .A(\u0_ps2_kb/_0107_ ), .Z(\u0_ps2_kb/_0011_ ) );
BUF_X1 \u0_ps2_kb/_1020_ ( .A(\u0_ps2_kb/_0090_ ), .Z(\u0_ps2_kb/_0186_ ) );
BUF_X1 \u0_ps2_kb/_1021_ ( .A(\u0_ps2_kb/_0108_ ), .Z(\u0_ps2_kb/_0012_ ) );
BUF_X1 \u0_ps2_kb/_1022_ ( .A(\u0_ps2_kb/_0091_ ), .Z(\u0_ps2_kb/_0187_ ) );
BUF_X1 \u0_ps2_kb/_1023_ ( .A(\u0_ps2_kb/_0109_ ), .Z(\u0_ps2_kb/_0013_ ) );
BUF_X1 \u0_ps2_kb/_1024_ ( .A(nextdata_n ), .Z(\u0_ps2_kb/_0471_ ) );
BUF_X1 \u0_ps2_kb/_1025_ ( .A(\u0_ps2_kb/_0092_ ), .Z(\u0_ps2_kb/_0188_ ) );
BUF_X1 \u0_ps2_kb/_1026_ ( .A(ready ), .Z(\u0_ps2_kb/_0479_ ) );
BUF_X1 \u0_ps2_kb/_1027_ ( .A(\u0_ps2_kb/_0111_ ), .Z(\u0_ps2_kb/_0015_ ) );
BUF_X1 \u0_ps2_kb/_1028_ ( .A(\u0_ps2_kb/_0087_ ), .Z(\u0_ps2_kb/_0183_ ) );
BUF_X1 \u0_ps2_kb/_1029_ ( .A(\u0_ps2_kb/_0112_ ), .Z(\u0_ps2_kb/_0016_ ) );
BUF_X1 \u0_ps2_kb/_1030_ ( .A(\u0_ps2_kb/_0086_ ), .Z(\u0_ps2_kb/_0182_ ) );
BUF_X1 \u0_ps2_kb/_1031_ ( .A(\u0_ps2_kb/_0113_ ), .Z(\u0_ps2_kb/_0017_ ) );
BUF_X1 \u0_ps2_kb/_1032_ ( .A(\u0_ps2_kb/_0115_ ), .Z(\u0_ps2_kb/_0019_ ) );
BUF_X1 \u0_ps2_kb/_1033_ ( .A(\u0_ps2_kb/_0093_ ), .Z(\u0_ps2_kb/_0189_ ) );
BUF_X1 \u0_ps2_kb/_1034_ ( .A(\u0_ps2_kb/_0116_ ), .Z(\u0_ps2_kb/_0020_ ) );
BUF_X1 \u0_ps2_kb/_1035_ ( .A(\u0_ps2_kb/_0094_ ), .Z(\u0_ps2_kb/_0190_ ) );
BUF_X1 \u0_ps2_kb/_1036_ ( .A(\u0_ps2_kb/_0117_ ), .Z(\u0_ps2_kb/_0021_ ) );
BUF_X1 \u0_ps2_kb/_1037_ ( .A(\u0_ps2_kb/_0104_ ), .Z(\u0_ps2_kb/_0008_ ) );
BUF_X1 \u0_ps2_kb/_1038_ ( .A(\u0_ps2_kb/_0105_ ), .Z(\u0_ps2_kb/_0009_ ) );
BUF_X1 \u0_ps2_kb/_1039_ ( .A(\u0_ps2_kb/_0114_ ), .Z(\u0_ps2_kb/_0018_ ) );
BUF_X1 \u0_ps2_kb/_1040_ ( .A(overflow ), .Z(\u0_ps2_kb/_0472_ ) );
BUF_X1 \u0_ps2_kb/_1041_ ( .A(\u0_ps2_kb/_0095_ ), .Z(\u0_ps2_kb/_0191_ ) );
BUF_X1 \u0_ps2_kb/_1042_ ( .A(\u0_ps2_kb/_0110_ ), .Z(\u0_ps2_kb/_0014_ ) );
DFF_X1 \u0_ps2_kb/_1043_ ( .D(\u0_ps2_kb/_0015_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr[0] ), .QN(\u0_ps2_kb/_0092_ ) );
DFF_X1 \u0_ps2_kb/_1044_ ( .D(\u0_ps2_kb/_0016_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr[1] ), .QN(\u0_ps2_kb/_0087_ ) );
DFF_X1 \u0_ps2_kb/_1045_ ( .D(\u0_ps2_kb/_0017_ ), .CK(clk ), .Q(\u0_ps2_kb/r_ptr[2] ), .QN(\u0_ps2_kb/_0086_ ) );
DFF_X1 \u0_ps2_kb/_1046_ ( .D(\u0_ps2_kb/_0078_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][0] ), .QN(\u0_ps2_kb/_0483_ ) );
DFF_X1 \u0_ps2_kb/_1047_ ( .D(\u0_ps2_kb/_0079_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][1] ), .QN(\u0_ps2_kb/_0484_ ) );
DFF_X1 \u0_ps2_kb/_1048_ ( .D(\u0_ps2_kb/_0080_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][2] ), .QN(\u0_ps2_kb/_0485_ ) );
DFF_X1 \u0_ps2_kb/_1049_ ( .D(\u0_ps2_kb/_0081_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][3] ), .QN(\u0_ps2_kb/_0486_ ) );
DFF_X1 \u0_ps2_kb/_1050_ ( .D(\u0_ps2_kb/_0082_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][4] ), .QN(\u0_ps2_kb/_0487_ ) );
DFF_X1 \u0_ps2_kb/_1051_ ( .D(\u0_ps2_kb/_0083_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][5] ), .QN(\u0_ps2_kb/_0488_ ) );
DFF_X1 \u0_ps2_kb/_1052_ ( .D(\u0_ps2_kb/_0084_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][6] ), .QN(\u0_ps2_kb/_0489_ ) );
DFF_X1 \u0_ps2_kb/_1053_ ( .D(\u0_ps2_kb/_0085_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[7][7] ), .QN(\u0_ps2_kb/_0490_ ) );
DFF_X1 \u0_ps2_kb/_1054_ ( .D(\u0_ps2_kb/_0070_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][0] ), .QN(\u0_ps2_kb/_0491_ ) );
DFF_X1 \u0_ps2_kb/_1055_ ( .D(\u0_ps2_kb/_0071_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][1] ), .QN(\u0_ps2_kb/_0492_ ) );
DFF_X1 \u0_ps2_kb/_1056_ ( .D(\u0_ps2_kb/_0072_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][2] ), .QN(\u0_ps2_kb/_0493_ ) );
DFF_X1 \u0_ps2_kb/_1057_ ( .D(\u0_ps2_kb/_0073_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][3] ), .QN(\u0_ps2_kb/_0494_ ) );
DFF_X1 \u0_ps2_kb/_1058_ ( .D(\u0_ps2_kb/_0074_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][4] ), .QN(\u0_ps2_kb/_0495_ ) );
DFF_X1 \u0_ps2_kb/_1059_ ( .D(\u0_ps2_kb/_0075_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][5] ), .QN(\u0_ps2_kb/_0496_ ) );
DFF_X1 \u0_ps2_kb/_1060_ ( .D(\u0_ps2_kb/_0076_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][6] ), .QN(\u0_ps2_kb/_0497_ ) );
DFF_X1 \u0_ps2_kb/_1061_ ( .D(\u0_ps2_kb/_0077_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[6][7] ), .QN(\u0_ps2_kb/_0498_ ) );
DFF_X1 \u0_ps2_kb/_1062_ ( .D(\u0_ps2_kb/_0062_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][0] ), .QN(\u0_ps2_kb/_0499_ ) );
DFF_X1 \u0_ps2_kb/_1063_ ( .D(\u0_ps2_kb/_0063_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][1] ), .QN(\u0_ps2_kb/_0500_ ) );
DFF_X1 \u0_ps2_kb/_1064_ ( .D(\u0_ps2_kb/_0064_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][2] ), .QN(\u0_ps2_kb/_0501_ ) );
DFF_X1 \u0_ps2_kb/_1065_ ( .D(\u0_ps2_kb/_0065_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][3] ), .QN(\u0_ps2_kb/_0502_ ) );
DFF_X1 \u0_ps2_kb/_1066_ ( .D(\u0_ps2_kb/_0066_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][4] ), .QN(\u0_ps2_kb/_0503_ ) );
DFF_X1 \u0_ps2_kb/_1067_ ( .D(\u0_ps2_kb/_0067_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][5] ), .QN(\u0_ps2_kb/_0504_ ) );
DFF_X1 \u0_ps2_kb/_1068_ ( .D(\u0_ps2_kb/_0068_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][6] ), .QN(\u0_ps2_kb/_0505_ ) );
DFF_X1 \u0_ps2_kb/_1069_ ( .D(\u0_ps2_kb/_0069_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[5][7] ), .QN(\u0_ps2_kb/_0506_ ) );
DFF_X1 \u0_ps2_kb/_1070_ ( .D(\u0_ps2_kb/_0054_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][0] ), .QN(\u0_ps2_kb/_0507_ ) );
DFF_X1 \u0_ps2_kb/_1071_ ( .D(\u0_ps2_kb/_0055_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][1] ), .QN(\u0_ps2_kb/_0508_ ) );
DFF_X1 \u0_ps2_kb/_1072_ ( .D(\u0_ps2_kb/_0056_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][2] ), .QN(\u0_ps2_kb/_0509_ ) );
DFF_X1 \u0_ps2_kb/_1073_ ( .D(\u0_ps2_kb/_0057_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][3] ), .QN(\u0_ps2_kb/_0510_ ) );
DFF_X1 \u0_ps2_kb/_1074_ ( .D(\u0_ps2_kb/_0058_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][4] ), .QN(\u0_ps2_kb/_0511_ ) );
DFF_X1 \u0_ps2_kb/_1075_ ( .D(\u0_ps2_kb/_0059_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][5] ), .QN(\u0_ps2_kb/_0512_ ) );
DFF_X1 \u0_ps2_kb/_1076_ ( .D(\u0_ps2_kb/_0060_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][6] ), .QN(\u0_ps2_kb/_0513_ ) );
DFF_X1 \u0_ps2_kb/_1077_ ( .D(\u0_ps2_kb/_0061_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[4][7] ), .QN(\u0_ps2_kb/_0514_ ) );
DFF_X1 \u0_ps2_kb/_1078_ ( .D(\u0_ps2_kb/_0038_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][0] ), .QN(\u0_ps2_kb/_0515_ ) );
DFF_X1 \u0_ps2_kb/_1079_ ( .D(\u0_ps2_kb/_0039_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][1] ), .QN(\u0_ps2_kb/_0516_ ) );
DFF_X1 \u0_ps2_kb/_1080_ ( .D(\u0_ps2_kb/_0040_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][2] ), .QN(\u0_ps2_kb/_0517_ ) );
DFF_X1 \u0_ps2_kb/_1081_ ( .D(\u0_ps2_kb/_0041_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][3] ), .QN(\u0_ps2_kb/_0518_ ) );
DFF_X1 \u0_ps2_kb/_1082_ ( .D(\u0_ps2_kb/_0042_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][4] ), .QN(\u0_ps2_kb/_0519_ ) );
DFF_X1 \u0_ps2_kb/_1083_ ( .D(\u0_ps2_kb/_0043_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][5] ), .QN(\u0_ps2_kb/_0520_ ) );
DFF_X1 \u0_ps2_kb/_1084_ ( .D(\u0_ps2_kb/_0044_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][6] ), .QN(\u0_ps2_kb/_0521_ ) );
DFF_X1 \u0_ps2_kb/_1085_ ( .D(\u0_ps2_kb/_0045_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[2][7] ), .QN(\u0_ps2_kb/_0522_ ) );
DFF_X1 \u0_ps2_kb/_1086_ ( .D(\u0_ps2_kb/_0046_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][0] ), .QN(\u0_ps2_kb/_0523_ ) );
DFF_X1 \u0_ps2_kb/_1087_ ( .D(\u0_ps2_kb/_0047_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][1] ), .QN(\u0_ps2_kb/_0524_ ) );
DFF_X1 \u0_ps2_kb/_1088_ ( .D(\u0_ps2_kb/_0048_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][2] ), .QN(\u0_ps2_kb/_0525_ ) );
DFF_X1 \u0_ps2_kb/_1089_ ( .D(\u0_ps2_kb/_0049_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][3] ), .QN(\u0_ps2_kb/_0526_ ) );
DFF_X1 \u0_ps2_kb/_1090_ ( .D(\u0_ps2_kb/_0050_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][4] ), .QN(\u0_ps2_kb/_0527_ ) );
DFF_X1 \u0_ps2_kb/_1091_ ( .D(\u0_ps2_kb/_0051_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][5] ), .QN(\u0_ps2_kb/_0528_ ) );
DFF_X1 \u0_ps2_kb/_1092_ ( .D(\u0_ps2_kb/_0052_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][6] ), .QN(\u0_ps2_kb/_0529_ ) );
DFF_X1 \u0_ps2_kb/_1093_ ( .D(\u0_ps2_kb/_0053_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[3][7] ), .QN(\u0_ps2_kb/_0530_ ) );
DFF_X1 \u0_ps2_kb/_1094_ ( .D(\u0_ps2_kb/_0022_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][0] ), .QN(\u0_ps2_kb/_0531_ ) );
DFF_X1 \u0_ps2_kb/_1095_ ( .D(\u0_ps2_kb/_0023_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][1] ), .QN(\u0_ps2_kb/_0532_ ) );
DFF_X1 \u0_ps2_kb/_1096_ ( .D(\u0_ps2_kb/_0024_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][2] ), .QN(\u0_ps2_kb/_0533_ ) );
DFF_X1 \u0_ps2_kb/_1097_ ( .D(\u0_ps2_kb/_0025_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][3] ), .QN(\u0_ps2_kb/_0534_ ) );
DFF_X1 \u0_ps2_kb/_1098_ ( .D(\u0_ps2_kb/_0026_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][4] ), .QN(\u0_ps2_kb/_0535_ ) );
DFF_X1 \u0_ps2_kb/_1099_ ( .D(\u0_ps2_kb/_0027_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][5] ), .QN(\u0_ps2_kb/_0536_ ) );
DFF_X1 \u0_ps2_kb/_1100_ ( .D(\u0_ps2_kb/_0028_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][6] ), .QN(\u0_ps2_kb/_0537_ ) );
DFF_X1 \u0_ps2_kb/_1101_ ( .D(\u0_ps2_kb/_0029_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[0][7] ), .QN(\u0_ps2_kb/_0538_ ) );
DFF_X1 \u0_ps2_kb/_1102_ ( .D(\u0_ps2_kb/_0030_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][0] ), .QN(\u0_ps2_kb/_0539_ ) );
DFF_X1 \u0_ps2_kb/_1103_ ( .D(\u0_ps2_kb/_0031_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][1] ), .QN(\u0_ps2_kb/_0540_ ) );
DFF_X1 \u0_ps2_kb/_1104_ ( .D(\u0_ps2_kb/_0032_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][2] ), .QN(\u0_ps2_kb/_0541_ ) );
DFF_X1 \u0_ps2_kb/_1105_ ( .D(\u0_ps2_kb/_0033_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][3] ), .QN(\u0_ps2_kb/_0542_ ) );
DFF_X1 \u0_ps2_kb/_1106_ ( .D(\u0_ps2_kb/_0034_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][4] ), .QN(\u0_ps2_kb/_0543_ ) );
DFF_X1 \u0_ps2_kb/_1107_ ( .D(\u0_ps2_kb/_0035_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][5] ), .QN(\u0_ps2_kb/_0544_ ) );
DFF_X1 \u0_ps2_kb/_1108_ ( .D(\u0_ps2_kb/_0036_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][6] ), .QN(\u0_ps2_kb/_0545_ ) );
DFF_X1 \u0_ps2_kb/_1109_ ( .D(\u0_ps2_kb/_0037_ ), .CK(clk ), .Q(\u0_ps2_kb/fifo[1][7] ), .QN(\u0_ps2_kb/_0546_ ) );
DFF_X1 \u0_ps2_kb/_1110_ ( .D(\u0_ps2_kb/_0014_ ), .CK(clk ), .Q(overflow ), .QN(\u0_ps2_kb/_0095_ ) );
DFF_X1 \u0_ps2_kb/_1111_ ( .D(\u0_ps2_kb/_0018_ ), .CK(clk ), .Q(ready ), .QN(\u0_ps2_kb/_0547_ ) );
DFF_X1 \u0_ps2_kb/_1112_ ( .D(\u0_ps2_kb/_0000_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[0] ), .QN(\u0_ps2_kb/_0548_ ) );
DFF_X1 \u0_ps2_kb/_1113_ ( .D(\u0_ps2_kb/_0001_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[1] ), .QN(\u0_ps2_kb/_0549_ ) );
DFF_X1 \u0_ps2_kb/_1114_ ( .D(\u0_ps2_kb/_0002_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[2] ), .QN(\u0_ps2_kb/_0550_ ) );
DFF_X1 \u0_ps2_kb/_1115_ ( .D(\u0_ps2_kb/_0003_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[3] ), .QN(\u0_ps2_kb/_0551_ ) );
DFF_X1 \u0_ps2_kb/_1116_ ( .D(\u0_ps2_kb/_0004_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[4] ), .QN(\u0_ps2_kb/_0552_ ) );
DFF_X1 \u0_ps2_kb/_1117_ ( .D(\u0_ps2_kb/_0005_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[5] ), .QN(\u0_ps2_kb/_0553_ ) );
DFF_X1 \u0_ps2_kb/_1118_ ( .D(\u0_ps2_kb/_0006_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[6] ), .QN(\u0_ps2_kb/_0554_ ) );
DFF_X1 \u0_ps2_kb/_1119_ ( .D(\u0_ps2_kb/_0007_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[7] ), .QN(\u0_ps2_kb/_0555_ ) );
DFF_X1 \u0_ps2_kb/_1120_ ( .D(\u0_ps2_kb/_0008_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[8] ), .QN(\u0_ps2_kb/_0556_ ) );
DFF_X1 \u0_ps2_kb/_1121_ ( .D(\u0_ps2_kb/_0009_ ), .CK(clk ), .Q(\u0_ps2_kb/buffer[9] ), .QN(\u0_ps2_kb/_0557_ ) );
DFF_X1 \u0_ps2_kb/_1122_ ( .D(\u0_ps2_kb/_0019_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr[0] ), .QN(\u0_ps2_kb/_0088_ ) );
DFF_X1 \u0_ps2_kb/_1123_ ( .D(\u0_ps2_kb/_0020_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr[1] ), .QN(\u0_ps2_kb/_0093_ ) );
DFF_X1 \u0_ps2_kb/_1124_ ( .D(\u0_ps2_kb/_0021_ ), .CK(clk ), .Q(\u0_ps2_kb/w_ptr[2] ), .QN(\u0_ps2_kb/_0094_ ) );
DFF_X1 \u0_ps2_kb/_1125_ ( .D(\u0_ps2_kb/_0010_ ), .CK(clk ), .Q(\u0_ps2_kb/count[0] ), .QN(\u0_ps2_kb/_0558_ ) );
DFF_X1 \u0_ps2_kb/_1126_ ( .D(\u0_ps2_kb/_0011_ ), .CK(clk ), .Q(\u0_ps2_kb/count[1] ), .QN(\u0_ps2_kb/_0089_ ) );
DFF_X1 \u0_ps2_kb/_1127_ ( .D(\u0_ps2_kb/_0012_ ), .CK(clk ), .Q(\u0_ps2_kb/count[2] ), .QN(\u0_ps2_kb/_0090_ ) );
DFF_X1 \u0_ps2_kb/_1128_ ( .D(\u0_ps2_kb/_0013_ ), .CK(clk ), .Q(\u0_ps2_kb/count[3] ), .QN(\u0_ps2_kb/_0091_ ) );
DFF_X1 \u0_ps2_kb/_1129_ ( .D(ps2_clk ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync[0] ), .QN(\u0_ps2_kb/_0559_ ) );
DFF_X1 \u0_ps2_kb/_1130_ ( .D(\u0_ps2_kb/ps2_clk_sync[0] ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync[1] ), .QN(\u0_ps2_kb/_0560_ ) );
DFF_X1 \u0_ps2_kb/_1131_ ( .D(\u0_ps2_kb/ps2_clk_sync[1] ), .CK(clk ), .Q(\u0_ps2_kb/ps2_clk_sync[2] ), .QN(\u0_ps2_kb/_0561_ ) );
NOR4_X2 \u1_ps2_dsh/_052_ ( .A1(\u1_ps2_dsh/_027_ ), .A2(\u1_ps2_dsh/_026_ ), .A3(\u1_ps2_dsh/_029_ ), .A4(\u1_ps2_dsh/_028_ ), .ZN(\u1_ps2_dsh/_034_ ) );
AND4_X1 \u1_ps2_dsh/_053_ ( .A1(\u1_ps2_dsh/_031_ ), .A2(\u1_ps2_dsh/_030_ ), .A3(\u1_ps2_dsh/_033_ ), .A4(\u1_ps2_dsh/_032_ ), .ZN(\u1_ps2_dsh/_035_ ) );
AND2_X1 \u1_ps2_dsh/_054_ ( .A1(\u1_ps2_dsh/_034_ ), .A2(\u1_ps2_dsh/_035_ ), .ZN(\u1_ps2_dsh/_017_ ) );
NAND2_X1 \u1_ps2_dsh/_055_ ( .A1(\u1_ps2_dsh/_031_ ), .A2(\u1_ps2_dsh/_032_ ), .ZN(\u1_ps2_dsh/_036_ ) );
NOR3_X2 \u1_ps2_dsh/_056_ ( .A1(\u1_ps2_dsh/_036_ ), .A2(\u1_ps2_dsh/_026_ ), .A3(\u1_ps2_dsh/_029_ ), .ZN(\u1_ps2_dsh/_037_ ) );
NAND2_X1 \u1_ps2_dsh/_057_ ( .A1(\u1_ps2_dsh/_030_ ), .A2(\u1_ps2_dsh/_033_ ), .ZN(\u1_ps2_dsh/_038_ ) );
NOR3_X2 \u1_ps2_dsh/_058_ ( .A1(\u1_ps2_dsh/_038_ ), .A2(\u1_ps2_dsh/_027_ ), .A3(\u1_ps2_dsh/_028_ ), .ZN(\u1_ps2_dsh/_039_ ) );
NAND2_X2 \u1_ps2_dsh/_059_ ( .A1(\u1_ps2_dsh/_037_ ), .A2(\u1_ps2_dsh/_039_ ), .ZN(\u1_ps2_dsh/_040_ ) );
AND2_X1 \u1_ps2_dsh/_060_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_018_ ), .ZN(\u1_ps2_dsh/_009_ ) );
AND2_X1 \u1_ps2_dsh/_061_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_019_ ), .ZN(\u1_ps2_dsh/_010_ ) );
AND2_X1 \u1_ps2_dsh/_062_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_020_ ), .ZN(\u1_ps2_dsh/_011_ ) );
AND2_X1 \u1_ps2_dsh/_063_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_021_ ), .ZN(\u1_ps2_dsh/_012_ ) );
AND2_X1 \u1_ps2_dsh/_064_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_022_ ), .ZN(\u1_ps2_dsh/_013_ ) );
AND2_X1 \u1_ps2_dsh/_065_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_023_ ), .ZN(\u1_ps2_dsh/_014_ ) );
AND2_X1 \u1_ps2_dsh/_066_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_024_ ), .ZN(\u1_ps2_dsh/_015_ ) );
AND2_X1 \u1_ps2_dsh/_067_ ( .A1(\u1_ps2_dsh/_040_ ), .A2(\u1_ps2_dsh/_025_ ), .ZN(\u1_ps2_dsh/_016_ ) );
LOGIC1_X1 \u1_ps2_dsh/_068_ ( .Z(\u1_ps2_dsh/_050_ ) );
LOGIC0_X1 \u1_ps2_dsh/_069_ ( .Z(\u1_ps2_dsh/_051_ ) );
BUF_X1 \u1_ps2_dsh/_070_ ( .A(\data_d1[1] ), .Z(\u1_ps2_dsh/_027_ ) );
BUF_X1 \u1_ps2_dsh/_071_ ( .A(\data_d1[0] ), .Z(\u1_ps2_dsh/_026_ ) );
BUF_X1 \u1_ps2_dsh/_072_ ( .A(\data_d1[3] ), .Z(\u1_ps2_dsh/_029_ ) );
BUF_X1 \u1_ps2_dsh/_073_ ( .A(\data_d1[2] ), .Z(\u1_ps2_dsh/_028_ ) );
BUF_X1 \u1_ps2_dsh/_074_ ( .A(\data_d1[5] ), .Z(\u1_ps2_dsh/_031_ ) );
BUF_X1 \u1_ps2_dsh/_075_ ( .A(\data_d1[4] ), .Z(\u1_ps2_dsh/_030_ ) );
BUF_X1 \u1_ps2_dsh/_076_ ( .A(\data_d1[7] ), .Z(\u1_ps2_dsh/_033_ ) );
BUF_X1 \u1_ps2_dsh/_077_ ( .A(\data_d1[6] ), .Z(\u1_ps2_dsh/_032_ ) );
BUF_X1 \u1_ps2_dsh/_078_ ( .A(\u1_ps2_dsh/_017_ ), .Z(\u1_ps2_dsh/_008_ ) );
BUF_X1 \u1_ps2_dsh/_079_ ( .A(\u1_ps2_dsh/ascii_result[0] ), .Z(\u1_ps2_dsh/_018_ ) );
BUF_X1 \u1_ps2_dsh/_080_ ( .A(\u1_ps2_dsh/_009_ ), .Z(\u1_ps2_dsh/_000_ ) );
BUF_X1 \u1_ps2_dsh/_081_ ( .A(\u1_ps2_dsh/ascii_result[1] ), .Z(\u1_ps2_dsh/_019_ ) );
BUF_X1 \u1_ps2_dsh/_082_ ( .A(\u1_ps2_dsh/_010_ ), .Z(\u1_ps2_dsh/_001_ ) );
BUF_X1 \u1_ps2_dsh/_083_ ( .A(\u1_ps2_dsh/ascii_result[2] ), .Z(\u1_ps2_dsh/_020_ ) );
BUF_X1 \u1_ps2_dsh/_084_ ( .A(\u1_ps2_dsh/_011_ ), .Z(\u1_ps2_dsh/_002_ ) );
BUF_X1 \u1_ps2_dsh/_085_ ( .A(\u1_ps2_dsh/ascii_result[3] ), .Z(\u1_ps2_dsh/_021_ ) );
BUF_X1 \u1_ps2_dsh/_086_ ( .A(\u1_ps2_dsh/_012_ ), .Z(\u1_ps2_dsh/_003_ ) );
BUF_X1 \u1_ps2_dsh/_087_ ( .A(\u1_ps2_dsh/ascii_result[4] ), .Z(\u1_ps2_dsh/_022_ ) );
BUF_X1 \u1_ps2_dsh/_088_ ( .A(\u1_ps2_dsh/_013_ ), .Z(\u1_ps2_dsh/_004_ ) );
BUF_X1 \u1_ps2_dsh/_089_ ( .A(\u1_ps2_dsh/ascii_result[5] ), .Z(\u1_ps2_dsh/_023_ ) );
BUF_X1 \u1_ps2_dsh/_090_ ( .A(\u1_ps2_dsh/_014_ ), .Z(\u1_ps2_dsh/_005_ ) );
BUF_X1 \u1_ps2_dsh/_091_ ( .A(\u1_ps2_dsh/ascii_result[6] ), .Z(\u1_ps2_dsh/_024_ ) );
BUF_X1 \u1_ps2_dsh/_092_ ( .A(\u1_ps2_dsh/_015_ ), .Z(\u1_ps2_dsh/_006_ ) );
BUF_X1 \u1_ps2_dsh/_093_ ( .A(\u1_ps2_dsh/ascii_result[7] ), .Z(\u1_ps2_dsh/_025_ ) );
BUF_X1 \u1_ps2_dsh/_094_ ( .A(\u1_ps2_dsh/_016_ ), .Z(\u1_ps2_dsh/_007_ ) );
DFFR_X1 \u1_ps2_dsh/_095_ ( .D(\u1_ps2_dsh/_008_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(key_release ), .QN(\u1_ps2_dsh/_041_ ) );
DFFR_X1 \u1_ps2_dsh/_096_ ( .D(\u1_ps2_dsh/_000_ ), .RN(fanout_net_2 ), .CK(clk ), .Q(\ascii[0] ), .QN(\u1_ps2_dsh/_042_ ) );
DFFR_X1 \u1_ps2_dsh/_097_ ( .D(\u1_ps2_dsh/_001_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[1] ), .QN(\u1_ps2_dsh/_043_ ) );
DFFR_X1 \u1_ps2_dsh/_098_ ( .D(\u1_ps2_dsh/_002_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[2] ), .QN(\u1_ps2_dsh/_044_ ) );
DFFR_X1 \u1_ps2_dsh/_099_ ( .D(\u1_ps2_dsh/_003_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[3] ), .QN(\u1_ps2_dsh/_045_ ) );
DFFR_X1 \u1_ps2_dsh/_100_ ( .D(\u1_ps2_dsh/_004_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[4] ), .QN(\u1_ps2_dsh/_046_ ) );
DFFR_X1 \u1_ps2_dsh/_101_ ( .D(\u1_ps2_dsh/_005_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[5] ), .QN(\u1_ps2_dsh/_047_ ) );
DFFR_X1 \u1_ps2_dsh/_102_ ( .D(\u1_ps2_dsh/_006_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[6] ), .QN(\u1_ps2_dsh/_048_ ) );
DFFR_X1 \u1_ps2_dsh/_103_ ( .D(\u1_ps2_dsh/_007_ ), .RN(clrn ), .CK(clk ), .Q(\ascii[7] ), .QN(\u1_ps2_dsh/_049_ ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_0_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[0] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_1_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[1] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_2_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[2] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_3_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[3] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_4_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[4] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_5_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[5] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_6_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[6] ) );
BUF_X1 \u1_ps2_dsh/key_ascii/i0/_7_ ( .A(\u1_ps2_dsh/_051_ ), .Z(\u1_ps2_dsh/ascii_result[7] ) );
INV_X32 \u2_ps2_cer/_067_ ( .A(\u2_ps2_cer/_056_ ), .ZN(\u2_ps2_cer/_021_ ) );
AND2_X4 \u2_ps2_cer/_068_ ( .A1(\u2_ps2_cer/_021_ ), .A2(\u2_ps2_cer/_057_ ), .ZN(\u2_ps2_cer/_022_ ) );
INV_X32 \u2_ps2_cer/_069_ ( .A(\u2_ps2_cer/_054_ ), .ZN(\u2_ps2_cer/_023_ ) );
NOR2_X4 \u2_ps2_cer/_070_ ( .A1(\u2_ps2_cer/_023_ ), .A2(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_024_ ) );
AND2_X4 \u2_ps2_cer/_071_ ( .A1(\u2_ps2_cer/_022_ ), .A2(\u2_ps2_cer/_024_ ), .ZN(\u2_ps2_cer/_025_ ) );
INV_X32 \u2_ps2_cer/_072_ ( .A(\u2_ps2_cer/_018_ ), .ZN(\u2_ps2_cer/_026_ ) );
AND2_X4 \u2_ps2_cer/_073_ ( .A1(\u2_ps2_cer/_026_ ), .A2(\u2_ps2_cer/_019_ ), .ZN(\u2_ps2_cer/_027_ ) );
AND2_X4 \u2_ps2_cer/_074_ ( .A1(\u2_ps2_cer/_025_ ), .A2(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_028_ ) );
INV_X16 \u2_ps2_cer/_075_ ( .A(\u2_ps2_cer/_050_ ), .ZN(\u2_ps2_cer/_029_ ) );
XNOR2_X1 \u2_ps2_cer/_076_ ( .A(\u2_ps2_cer/_028_ ), .B(\u2_ps2_cer/_029_ ), .ZN(\u2_ps2_cer/_010_ ) );
NOR2_X1 \u2_ps2_cer/_077_ ( .A1(\u2_ps2_cer/_029_ ), .A2(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_030_ ) );
INV_X2 \u2_ps2_cer/_078_ ( .A(\u2_ps2_cer/_053_ ), .ZN(\u2_ps2_cer/_031_ ) );
OAI211_X2 \u2_ps2_cer/_079_ ( .A(\u2_ps2_cer/_028_ ), .B(\u2_ps2_cer/_030_ ), .C1(\u2_ps2_cer/_052_ ), .C2(\u2_ps2_cer/_031_ ), .ZN(\u2_ps2_cer/_032_ ) );
INV_X1 \u2_ps2_cer/_080_ ( .A(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_033_ ) );
AND3_X1 \u2_ps2_cer/_081_ ( .A1(\u2_ps2_cer/_025_ ), .A2(\u2_ps2_cer/_050_ ), .A3(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_034_ ) );
OAI21_X1 \u2_ps2_cer/_082_ ( .A(\u2_ps2_cer/_032_ ), .B1(\u2_ps2_cer/_033_ ), .B2(\u2_ps2_cer/_034_ ), .ZN(\u2_ps2_cer/_011_ ) );
AND2_X4 \u2_ps2_cer/_083_ ( .A1(\u2_ps2_cer/_050_ ), .A2(\u2_ps2_cer/_051_ ), .ZN(\u2_ps2_cer/_035_ ) );
NAND2_X2 \u2_ps2_cer/_084_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_035_ ), .ZN(\u2_ps2_cer/_036_ ) );
XNOR2_X1 \u2_ps2_cer/_085_ ( .A(\u2_ps2_cer/_036_ ), .B(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_012_ ) );
NAND4_X1 \u2_ps2_cer/_086_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_052_ ), .A3(\u2_ps2_cer/_031_ ), .A4(\u2_ps2_cer/_035_ ), .ZN(\u2_ps2_cer/_037_ ) );
INV_X1 \u2_ps2_cer/_087_ ( .A(\u2_ps2_cer/_028_ ), .ZN(\u2_ps2_cer/_038_ ) );
NOR2_X1 \u2_ps2_cer/_088_ ( .A1(\u2_ps2_cer/_031_ ), .A2(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_039_ ) );
AOI22_X1 \u2_ps2_cer/_089_ ( .A1(\u2_ps2_cer/_039_ ), .A2(\u2_ps2_cer/_030_ ), .B1(\u2_ps2_cer/_035_ ), .B2(\u2_ps2_cer/_052_ ), .ZN(\u2_ps2_cer/_040_ ) );
NOR2_X2 \u2_ps2_cer/_090_ ( .A1(\u2_ps2_cer/_038_ ), .A2(\u2_ps2_cer/_040_ ), .ZN(\u2_ps2_cer/_041_ ) );
OAI21_X1 \u2_ps2_cer/_091_ ( .A(\u2_ps2_cer/_037_ ), .B1(\u2_ps2_cer/_041_ ), .B2(\u2_ps2_cer/_031_ ), .ZN(\u2_ps2_cer/_013_ ) );
XNOR2_X1 \u2_ps2_cer/_092_ ( .A(\u2_ps2_cer/_027_ ), .B(\u2_ps2_cer/_023_ ), .ZN(\u2_ps2_cer/_014_ ) );
NAND3_X1 \u2_ps2_cer/_093_ ( .A1(\u2_ps2_cer/_024_ ), .A2(\u2_ps2_cer/_026_ ), .A3(\u2_ps2_cer/_019_ ), .ZN(\u2_ps2_cer/_042_ ) );
AND3_X4 \u2_ps2_cer/_094_ ( .A1(\u2_ps2_cer/_026_ ), .A2(\u2_ps2_cer/_019_ ), .A3(\u2_ps2_cer/_054_ ), .ZN(\u2_ps2_cer/_043_ ) );
INV_X1 \u2_ps2_cer/_095_ ( .A(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_044_ ) );
OAI22_X1 \u2_ps2_cer/_096_ ( .A1(\u2_ps2_cer/_042_ ), .A2(\u2_ps2_cer/_022_ ), .B1(\u2_ps2_cer/_043_ ), .B2(\u2_ps2_cer/_044_ ), .ZN(\u2_ps2_cer/_015_ ) );
AND2_X4 \u2_ps2_cer/_097_ ( .A1(\u2_ps2_cer/_054_ ), .A2(\u2_ps2_cer/_055_ ), .ZN(\u2_ps2_cer/_045_ ) );
AND2_X2 \u2_ps2_cer/_098_ ( .A1(\u2_ps2_cer/_027_ ), .A2(\u2_ps2_cer/_045_ ), .ZN(\u2_ps2_cer/_046_ ) );
XNOR2_X1 \u2_ps2_cer/_099_ ( .A(\u2_ps2_cer/_046_ ), .B(\u2_ps2_cer/_021_ ), .ZN(\u2_ps2_cer/_016_ ) );
AOI21_X1 \u2_ps2_cer/_100_ ( .A(\u2_ps2_cer/_057_ ), .B1(\u2_ps2_cer/_046_ ), .B2(\u2_ps2_cer/_056_ ), .ZN(\u2_ps2_cer/_047_ ) );
AND4_X1 \u2_ps2_cer/_101_ ( .A1(\u2_ps2_cer/_056_ ), .A2(\u2_ps2_cer/_027_ ), .A3(\u2_ps2_cer/_057_ ), .A4(\u2_ps2_cer/_045_ ), .ZN(\u2_ps2_cer/_048_ ) );
NOR3_X1 \u2_ps2_cer/_102_ ( .A1(\u2_ps2_cer/_028_ ), .A2(\u2_ps2_cer/_047_ ), .A3(\u2_ps2_cer/_048_ ), .ZN(\u2_ps2_cer/_017_ ) );
INV_X1 \u2_ps2_cer/_103_ ( .A(\u2_ps2_cer/_027_ ), .ZN(\u2_ps2_cer/_049_ ) );
OAI21_X1 \u2_ps2_cer/_104_ ( .A(\u2_ps2_cer/_049_ ), .B1(\u2_ps2_cer/_026_ ), .B2(\u2_ps2_cer/_020_ ), .ZN(\u2_ps2_cer/_009_ ) );
BUF_X1 \u2_ps2_cer/_105_ ( .A(\u2_ps2_cer/counted ), .Z(\u2_ps2_cer/_018_ ) );
BUF_X1 \u2_ps2_cer/_106_ ( .A(_026_ ), .Z(\u2_ps2_cer/_019_ ) );
BUF_X1 \u2_ps2_cer/_107_ ( .A(\high_tens[0] ), .Z(\u2_ps2_cer/_050_ ) );
BUF_X1 \u2_ps2_cer/_108_ ( .A(\high_tens[1] ), .Z(\u2_ps2_cer/_051_ ) );
BUF_X1 \u2_ps2_cer/_109_ ( .A(\high_tens[2] ), .Z(\u2_ps2_cer/_052_ ) );
BUF_X1 \u2_ps2_cer/_110_ ( .A(\high_tens[3] ), .Z(\u2_ps2_cer/_053_ ) );
BUF_X1 \u2_ps2_cer/_111_ ( .A(\high_units[0] ), .Z(\u2_ps2_cer/_054_ ) );
BUF_X1 \u2_ps2_cer/_112_ ( .A(\high_units[1] ), .Z(\u2_ps2_cer/_055_ ) );
BUF_X1 \u2_ps2_cer/_113_ ( .A(\high_units[2] ), .Z(\u2_ps2_cer/_056_ ) );
BUF_X1 \u2_ps2_cer/_114_ ( .A(\high_units[3] ), .Z(\u2_ps2_cer/_057_ ) );
BUF_X1 \u2_ps2_cer/_115_ ( .A(\u2_ps2_cer/_010_ ), .Z(\u2_ps2_cer/_001_ ) );
BUF_X1 \u2_ps2_cer/_116_ ( .A(\u2_ps2_cer/_011_ ), .Z(\u2_ps2_cer/_002_ ) );
BUF_X1 \u2_ps2_cer/_117_ ( .A(\u2_ps2_cer/_012_ ), .Z(\u2_ps2_cer/_003_ ) );
BUF_X1 \u2_ps2_cer/_118_ ( .A(\u2_ps2_cer/_013_ ), .Z(\u2_ps2_cer/_004_ ) );
BUF_X1 \u2_ps2_cer/_119_ ( .A(\u2_ps2_cer/_014_ ), .Z(\u2_ps2_cer/_005_ ) );
BUF_X1 \u2_ps2_cer/_120_ ( .A(\u2_ps2_cer/_015_ ), .Z(\u2_ps2_cer/_006_ ) );
BUF_X1 \u2_ps2_cer/_121_ ( .A(\u2_ps2_cer/_016_ ), .Z(\u2_ps2_cer/_007_ ) );
BUF_X1 \u2_ps2_cer/_122_ ( .A(\u2_ps2_cer/_017_ ), .Z(\u2_ps2_cer/_008_ ) );
BUF_X1 \u2_ps2_cer/_123_ ( .A(key_release ), .Z(\u2_ps2_cer/_020_ ) );
BUF_X1 \u2_ps2_cer/_124_ ( .A(\u2_ps2_cer/_009_ ), .Z(\u2_ps2_cer/_000_ ) );
DFFR_X1 \u2_ps2_cer/_125_ ( .D(\u2_ps2_cer/_005_ ), .RN(clrn ), .CK(clk ), .Q(\high_units[0] ), .QN(\u2_ps2_cer/_058_ ) );
DFFR_X1 \u2_ps2_cer/_126_ ( .D(\u2_ps2_cer/_006_ ), .RN(clrn ), .CK(clk ), .Q(\high_units[1] ), .QN(\u2_ps2_cer/_059_ ) );
DFFR_X1 \u2_ps2_cer/_127_ ( .D(\u2_ps2_cer/_007_ ), .RN(clrn ), .CK(clk ), .Q(\high_units[2] ), .QN(\u2_ps2_cer/_060_ ) );
DFFR_X1 \u2_ps2_cer/_128_ ( .D(\u2_ps2_cer/_008_ ), .RN(clrn ), .CK(clk ), .Q(\high_units[3] ), .QN(\u2_ps2_cer/_061_ ) );
DFFR_X1 \u2_ps2_cer/_129_ ( .D(\u2_ps2_cer/_001_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens[0] ), .QN(\u2_ps2_cer/_062_ ) );
DFFR_X1 \u2_ps2_cer/_130_ ( .D(\u2_ps2_cer/_002_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens[1] ), .QN(\u2_ps2_cer/_063_ ) );
DFFR_X1 \u2_ps2_cer/_131_ ( .D(\u2_ps2_cer/_003_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens[2] ), .QN(\u2_ps2_cer/_064_ ) );
DFFR_X1 \u2_ps2_cer/_132_ ( .D(\u2_ps2_cer/_004_ ), .RN(clrn ), .CK(clk ), .Q(\high_tens[3] ), .QN(\u2_ps2_cer/_065_ ) );
DFFR_X1 \u2_ps2_cer/_133_ ( .D(\u2_ps2_cer/_000_ ), .RN(clrn ), .CK(clk ), .Q(\u2_ps2_cer/counted ), .QN(\u2_ps2_cer/_066_ ) );
NOR2_X4 \u3_seg_h_0/_43_ ( .A1(\u3_seg_h_0/_31_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_01_ ) );
INV_X2 \u3_seg_h_0/_44_ ( .A(\u3_seg_h_0/_01_ ), .ZN(\u3_seg_h_0/_02_ ) );
INV_X4 \u3_seg_h_0/_45_ ( .A(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_03_ ) );
NOR2_X2 \u3_seg_h_0/_46_ ( .A1(\u3_seg_h_0/_03_ ), .A2(\u3_seg_h_0/_34_ ), .ZN(\u3_seg_h_0/_04_ ) );
INV_X16 \u3_seg_h_0/_47_ ( .A(\u3_seg_h_0/_34_ ), .ZN(\u3_seg_h_0/_05_ ) );
NOR2_X2 \u3_seg_h_0/_48_ ( .A1(\u3_seg_h_0/_05_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_06_ ) );
OR3_X4 \u3_seg_h_0/_49_ ( .A1(\u3_seg_h_0/_02_ ), .A2(\u3_seg_h_0/_04_ ), .A3(\u3_seg_h_0/_06_ ), .ZN(\u3_seg_h_0/_07_ ) );
INV_X32 \u3_seg_h_0/_50_ ( .A(\u3_seg_h_0/_31_ ), .ZN(\u3_seg_h_0/_08_ ) );
NOR2_X2 \u3_seg_h_0/_51_ ( .A1(\u3_seg_h_0/_08_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_09_ ) );
NOR2_X4 \u3_seg_h_0/_52_ ( .A1(\u3_seg_h_0/_34_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_10_ ) );
AND2_X1 \u3_seg_h_0/_53_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_10_ ), .ZN(\u3_seg_h_0/_11_ ) );
INV_X1 \u3_seg_h_0/_54_ ( .A(\u3_seg_h_0/_11_ ), .ZN(\u3_seg_h_0/_12_ ) );
INV_X1 \u3_seg_h_0/_55_ ( .A(\u3_seg_h_0/_00_ ), .ZN(\u3_seg_h_0/_13_ ) );
AND2_X4 \u3_seg_h_0/_56_ ( .A1(\u3_seg_h_0/_31_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_14_ ) );
AOI21_X1 \u3_seg_h_0/_57_ ( .A(\u3_seg_h_0/_13_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_15_ ) );
NAND3_X1 \u3_seg_h_0/_58_ ( .A1(\u3_seg_h_0/_07_ ), .A2(\u3_seg_h_0/_12_ ), .A3(\u3_seg_h_0/_15_ ), .ZN(\u3_seg_h_0/_35_ ) );
NAND2_X1 \u3_seg_h_0/_59_ ( .A1(\u3_seg_h_0/_02_ ), .A2(\u3_seg_h_0/_10_ ), .ZN(\u3_seg_h_0/_16_ ) );
AND2_X2 \u3_seg_h_0/_60_ ( .A1(\u3_seg_h_0/_34_ ), .A2(\u3_seg_h_0/_33_ ), .ZN(\u3_seg_h_0/_17_ ) );
NAND2_X1 \u3_seg_h_0/_61_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_17_ ), .ZN(\u3_seg_h_0/_18_ ) );
NAND3_X1 \u3_seg_h_0/_62_ ( .A1(\u3_seg_h_0/_15_ ), .A2(\u3_seg_h_0/_16_ ), .A3(\u3_seg_h_0/_18_ ), .ZN(\u3_seg_h_0/_36_ ) );
NOR3_X1 \u3_seg_h_0/_63_ ( .A1(\u3_seg_h_0/_03_ ), .A2(\u3_seg_h_0/_34_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_19_ ) );
AOI21_X1 \u3_seg_h_0/_64_ ( .A(\u3_seg_h_0/_19_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_20_ ) );
NAND3_X1 \u3_seg_h_0/_65_ ( .A1(\u3_seg_h_0/_05_ ), .A2(\u3_seg_h_0/_03_ ), .A3(\u3_seg_h_0/_31_ ), .ZN(\u3_seg_h_0/_21_ ) );
NAND2_X1 \u3_seg_h_0/_66_ ( .A1(\u3_seg_h_0/_09_ ), .A2(\u3_seg_h_0/_06_ ), .ZN(\u3_seg_h_0/_22_ ) );
NAND4_X1 \u3_seg_h_0/_67_ ( .A1(\u3_seg_h_0/_20_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_21_ ), .A4(\u3_seg_h_0/_22_ ), .ZN(\u3_seg_h_0/_37_ ) );
NAND3_X1 \u3_seg_h_0/_68_ ( .A1(\u3_seg_h_0/_06_ ), .A2(\u3_seg_h_0/_08_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_23_ ) );
AOI22_X1 \u3_seg_h_0/_69_ ( .A1(\u3_seg_h_0/_04_ ), .A2(\u3_seg_h_0/_01_ ), .B1(\u3_seg_h_0/_14_ ), .B2(\u3_seg_h_0/_17_ ), .ZN(\u3_seg_h_0/_24_ ) );
NAND4_X1 \u3_seg_h_0/_70_ ( .A1(\u3_seg_h_0/_12_ ), .A2(\u3_seg_h_0/_15_ ), .A3(\u3_seg_h_0/_23_ ), .A4(\u3_seg_h_0/_24_ ), .ZN(\u3_seg_h_0/_38_ ) );
OAI21_X1 \u3_seg_h_0/_71_ ( .A(\u3_seg_h_0/_17_ ), .B1(\u3_seg_h_0/_08_ ), .B2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_25_ ) );
NAND3_X1 \u3_seg_h_0/_72_ ( .A1(\u3_seg_h_0/_10_ ), .A2(\u3_seg_h_0/_08_ ), .A3(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_26_ ) );
NAND3_X1 \u3_seg_h_0/_73_ ( .A1(\u3_seg_h_0/_25_ ), .A2(\u3_seg_h_0/_26_ ), .A3(\u3_seg_h_0/_00_ ), .ZN(\u3_seg_h_0/_39_ ) );
AND2_X1 \u3_seg_h_0/_74_ ( .A1(\u3_seg_h_0/_08_ ), .A2(\u3_seg_h_0/_32_ ), .ZN(\u3_seg_h_0/_27_ ) );
OAI21_X1 \u3_seg_h_0/_75_ ( .A(\u3_seg_h_0/_04_ ), .B1(\u3_seg_h_0/_27_ ), .B2(\u3_seg_h_0/_09_ ), .ZN(\u3_seg_h_0/_28_ ) );
NAND2_X1 \u3_seg_h_0/_76_ ( .A1(\u3_seg_h_0/_06_ ), .A2(\u3_seg_h_0/_14_ ), .ZN(\u3_seg_h_0/_29_ ) );
NAND4_X1 \u3_seg_h_0/_77_ ( .A1(\u3_seg_h_0/_28_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_25_ ), .A4(\u3_seg_h_0/_29_ ), .ZN(\u3_seg_h_0/_40_ ) );
AOI22_X1 \u3_seg_h_0/_78_ ( .A1(\u3_seg_h_0/_10_ ), .A2(\u3_seg_h_0/_09_ ), .B1(\u3_seg_h_0/_04_ ), .B2(\u3_seg_h_0/_01_ ), .ZN(\u3_seg_h_0/_30_ ) );
NAND4_X1 \u3_seg_h_0/_79_ ( .A1(\u3_seg_h_0/_30_ ), .A2(\u3_seg_h_0/_00_ ), .A3(\u3_seg_h_0/_18_ ), .A4(\u3_seg_h_0/_29_ ), .ZN(\u3_seg_h_0/_41_ ) );
LOGIC1_X1 \u3_seg_h_0/_80_ ( .Z(\u3_seg_h_0/_42_ ) );
BUF_X1 \u3_seg_h_0/_81_ ( .A(\u3_seg_h_0/_42_ ), .Z(\seg_out_2[0] ) );
BUF_X1 \u3_seg_h_0/_82_ ( .A(\key_ascii_display[3] ), .Z(\u3_seg_h_0/_34_ ) );
BUF_X1 \u3_seg_h_0/_83_ ( .A(\key_ascii_display[2] ), .Z(\u3_seg_h_0/_33_ ) );
BUF_X1 \u3_seg_h_0/_84_ ( .A(\key_ascii_display[0] ), .Z(\u3_seg_h_0/_31_ ) );
BUF_X1 \u3_seg_h_0/_85_ ( .A(\key_ascii_display[1] ), .Z(\u3_seg_h_0/_32_ ) );
BUF_X1 \u3_seg_h_0/_86_ ( .A(en ), .Z(\u3_seg_h_0/_00_ ) );
BUF_X1 \u3_seg_h_0/_87_ ( .A(\u3_seg_h_0/_35_ ), .Z(\seg_out_2[1] ) );
BUF_X1 \u3_seg_h_0/_88_ ( .A(\u3_seg_h_0/_36_ ), .Z(\seg_out_2[2] ) );
BUF_X1 \u3_seg_h_0/_89_ ( .A(\u3_seg_h_0/_37_ ), .Z(\seg_out_2[3] ) );
BUF_X1 \u3_seg_h_0/_90_ ( .A(\u3_seg_h_0/_38_ ), .Z(\seg_out_2[4] ) );
BUF_X1 \u3_seg_h_0/_91_ ( .A(\u3_seg_h_0/_39_ ), .Z(\seg_out_2[5] ) );
BUF_X1 \u3_seg_h_0/_92_ ( .A(\u3_seg_h_0/_40_ ), .Z(\seg_out_2[6] ) );
BUF_X1 \u3_seg_h_0/_93_ ( .A(\u3_seg_h_0/_41_ ), .Z(\seg_out_2[7] ) );
NOR2_X4 \u4_seg_h_1/_43_ ( .A1(\u4_seg_h_1/_31_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_01_ ) );
INV_X2 \u4_seg_h_1/_44_ ( .A(\u4_seg_h_1/_01_ ), .ZN(\u4_seg_h_1/_02_ ) );
INV_X4 \u4_seg_h_1/_45_ ( .A(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_03_ ) );
NOR2_X2 \u4_seg_h_1/_46_ ( .A1(\u4_seg_h_1/_03_ ), .A2(\u4_seg_h_1/_34_ ), .ZN(\u4_seg_h_1/_04_ ) );
INV_X16 \u4_seg_h_1/_47_ ( .A(\u4_seg_h_1/_34_ ), .ZN(\u4_seg_h_1/_05_ ) );
NOR2_X2 \u4_seg_h_1/_48_ ( .A1(\u4_seg_h_1/_05_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_06_ ) );
OR3_X4 \u4_seg_h_1/_49_ ( .A1(\u4_seg_h_1/_02_ ), .A2(\u4_seg_h_1/_04_ ), .A3(\u4_seg_h_1/_06_ ), .ZN(\u4_seg_h_1/_07_ ) );
INV_X32 \u4_seg_h_1/_50_ ( .A(\u4_seg_h_1/_31_ ), .ZN(\u4_seg_h_1/_08_ ) );
NOR2_X2 \u4_seg_h_1/_51_ ( .A1(\u4_seg_h_1/_08_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_09_ ) );
NOR2_X4 \u4_seg_h_1/_52_ ( .A1(\u4_seg_h_1/_34_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_10_ ) );
AND2_X1 \u4_seg_h_1/_53_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_10_ ), .ZN(\u4_seg_h_1/_11_ ) );
INV_X1 \u4_seg_h_1/_54_ ( .A(\u4_seg_h_1/_11_ ), .ZN(\u4_seg_h_1/_12_ ) );
INV_X1 \u4_seg_h_1/_55_ ( .A(\u4_seg_h_1/_00_ ), .ZN(\u4_seg_h_1/_13_ ) );
AND2_X4 \u4_seg_h_1/_56_ ( .A1(\u4_seg_h_1/_31_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_14_ ) );
AOI21_X1 \u4_seg_h_1/_57_ ( .A(\u4_seg_h_1/_13_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_15_ ) );
NAND3_X1 \u4_seg_h_1/_58_ ( .A1(\u4_seg_h_1/_07_ ), .A2(\u4_seg_h_1/_12_ ), .A3(\u4_seg_h_1/_15_ ), .ZN(\u4_seg_h_1/_35_ ) );
NAND2_X1 \u4_seg_h_1/_59_ ( .A1(\u4_seg_h_1/_02_ ), .A2(\u4_seg_h_1/_10_ ), .ZN(\u4_seg_h_1/_16_ ) );
AND2_X2 \u4_seg_h_1/_60_ ( .A1(\u4_seg_h_1/_34_ ), .A2(\u4_seg_h_1/_33_ ), .ZN(\u4_seg_h_1/_17_ ) );
NAND2_X1 \u4_seg_h_1/_61_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_17_ ), .ZN(\u4_seg_h_1/_18_ ) );
NAND3_X1 \u4_seg_h_1/_62_ ( .A1(\u4_seg_h_1/_15_ ), .A2(\u4_seg_h_1/_16_ ), .A3(\u4_seg_h_1/_18_ ), .ZN(\u4_seg_h_1/_36_ ) );
NOR3_X1 \u4_seg_h_1/_63_ ( .A1(\u4_seg_h_1/_03_ ), .A2(\u4_seg_h_1/_34_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_19_ ) );
AOI21_X1 \u4_seg_h_1/_64_ ( .A(\u4_seg_h_1/_19_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_20_ ) );
NAND3_X1 \u4_seg_h_1/_65_ ( .A1(\u4_seg_h_1/_05_ ), .A2(\u4_seg_h_1/_03_ ), .A3(\u4_seg_h_1/_31_ ), .ZN(\u4_seg_h_1/_21_ ) );
NAND2_X1 \u4_seg_h_1/_66_ ( .A1(\u4_seg_h_1/_09_ ), .A2(\u4_seg_h_1/_06_ ), .ZN(\u4_seg_h_1/_22_ ) );
NAND4_X1 \u4_seg_h_1/_67_ ( .A1(\u4_seg_h_1/_20_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_21_ ), .A4(\u4_seg_h_1/_22_ ), .ZN(\u4_seg_h_1/_37_ ) );
NAND3_X1 \u4_seg_h_1/_68_ ( .A1(\u4_seg_h_1/_06_ ), .A2(\u4_seg_h_1/_08_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_23_ ) );
AOI22_X1 \u4_seg_h_1/_69_ ( .A1(\u4_seg_h_1/_04_ ), .A2(\u4_seg_h_1/_01_ ), .B1(\u4_seg_h_1/_14_ ), .B2(\u4_seg_h_1/_17_ ), .ZN(\u4_seg_h_1/_24_ ) );
NAND4_X1 \u4_seg_h_1/_70_ ( .A1(\u4_seg_h_1/_12_ ), .A2(\u4_seg_h_1/_15_ ), .A3(\u4_seg_h_1/_23_ ), .A4(\u4_seg_h_1/_24_ ), .ZN(\u4_seg_h_1/_38_ ) );
OAI21_X1 \u4_seg_h_1/_71_ ( .A(\u4_seg_h_1/_17_ ), .B1(\u4_seg_h_1/_08_ ), .B2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_25_ ) );
NAND3_X1 \u4_seg_h_1/_72_ ( .A1(\u4_seg_h_1/_10_ ), .A2(\u4_seg_h_1/_08_ ), .A3(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_26_ ) );
NAND3_X1 \u4_seg_h_1/_73_ ( .A1(\u4_seg_h_1/_25_ ), .A2(\u4_seg_h_1/_26_ ), .A3(\u4_seg_h_1/_00_ ), .ZN(\u4_seg_h_1/_39_ ) );
AND2_X1 \u4_seg_h_1/_74_ ( .A1(\u4_seg_h_1/_08_ ), .A2(\u4_seg_h_1/_32_ ), .ZN(\u4_seg_h_1/_27_ ) );
OAI21_X1 \u4_seg_h_1/_75_ ( .A(\u4_seg_h_1/_04_ ), .B1(\u4_seg_h_1/_27_ ), .B2(\u4_seg_h_1/_09_ ), .ZN(\u4_seg_h_1/_28_ ) );
NAND2_X1 \u4_seg_h_1/_76_ ( .A1(\u4_seg_h_1/_06_ ), .A2(\u4_seg_h_1/_14_ ), .ZN(\u4_seg_h_1/_29_ ) );
NAND4_X1 \u4_seg_h_1/_77_ ( .A1(\u4_seg_h_1/_28_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_25_ ), .A4(\u4_seg_h_1/_29_ ), .ZN(\u4_seg_h_1/_40_ ) );
AOI22_X1 \u4_seg_h_1/_78_ ( .A1(\u4_seg_h_1/_10_ ), .A2(\u4_seg_h_1/_09_ ), .B1(\u4_seg_h_1/_04_ ), .B2(\u4_seg_h_1/_01_ ), .ZN(\u4_seg_h_1/_30_ ) );
NAND4_X1 \u4_seg_h_1/_79_ ( .A1(\u4_seg_h_1/_30_ ), .A2(\u4_seg_h_1/_00_ ), .A3(\u4_seg_h_1/_18_ ), .A4(\u4_seg_h_1/_29_ ), .ZN(\u4_seg_h_1/_41_ ) );
LOGIC1_X1 \u4_seg_h_1/_80_ ( .Z(\u4_seg_h_1/_42_ ) );
BUF_X1 \u4_seg_h_1/_81_ ( .A(\u4_seg_h_1/_42_ ), .Z(\seg_out_3[0] ) );
BUF_X1 \u4_seg_h_1/_82_ ( .A(\key_ascii_display[7] ), .Z(\u4_seg_h_1/_34_ ) );
BUF_X1 \u4_seg_h_1/_83_ ( .A(\key_ascii_display[6] ), .Z(\u4_seg_h_1/_33_ ) );
BUF_X1 \u4_seg_h_1/_84_ ( .A(\key_ascii_display[4] ), .Z(\u4_seg_h_1/_31_ ) );
BUF_X1 \u4_seg_h_1/_85_ ( .A(\key_ascii_display[5] ), .Z(\u4_seg_h_1/_32_ ) );
BUF_X1 \u4_seg_h_1/_86_ ( .A(en ), .Z(\u4_seg_h_1/_00_ ) );
BUF_X1 \u4_seg_h_1/_87_ ( .A(\u4_seg_h_1/_35_ ), .Z(\seg_out_3[1] ) );
BUF_X1 \u4_seg_h_1/_88_ ( .A(\u4_seg_h_1/_36_ ), .Z(\seg_out_3[2] ) );
BUF_X1 \u4_seg_h_1/_89_ ( .A(\u4_seg_h_1/_37_ ), .Z(\seg_out_3[3] ) );
BUF_X1 \u4_seg_h_1/_90_ ( .A(\u4_seg_h_1/_38_ ), .Z(\seg_out_3[4] ) );
BUF_X1 \u4_seg_h_1/_91_ ( .A(\u4_seg_h_1/_39_ ), .Z(\seg_out_3[5] ) );
BUF_X1 \u4_seg_h_1/_92_ ( .A(\u4_seg_h_1/_40_ ), .Z(\seg_out_3[6] ) );
BUF_X1 \u4_seg_h_1/_93_ ( .A(\u4_seg_h_1/_41_ ), .Z(\seg_out_3[7] ) );
NOR2_X4 \u5_seg_h_2/_43_ ( .A1(\u5_seg_h_2/_31_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_01_ ) );
INV_X2 \u5_seg_h_2/_44_ ( .A(\u5_seg_h_2/_01_ ), .ZN(\u5_seg_h_2/_02_ ) );
INV_X4 \u5_seg_h_2/_45_ ( .A(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_03_ ) );
NOR2_X2 \u5_seg_h_2/_46_ ( .A1(\u5_seg_h_2/_03_ ), .A2(\u5_seg_h_2/_34_ ), .ZN(\u5_seg_h_2/_04_ ) );
INV_X16 \u5_seg_h_2/_47_ ( .A(\u5_seg_h_2/_34_ ), .ZN(\u5_seg_h_2/_05_ ) );
NOR2_X2 \u5_seg_h_2/_48_ ( .A1(\u5_seg_h_2/_05_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_06_ ) );
OR3_X4 \u5_seg_h_2/_49_ ( .A1(\u5_seg_h_2/_02_ ), .A2(\u5_seg_h_2/_04_ ), .A3(\u5_seg_h_2/_06_ ), .ZN(\u5_seg_h_2/_07_ ) );
INV_X32 \u5_seg_h_2/_50_ ( .A(\u5_seg_h_2/_31_ ), .ZN(\u5_seg_h_2/_08_ ) );
NOR2_X2 \u5_seg_h_2/_51_ ( .A1(\u5_seg_h_2/_08_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_09_ ) );
NOR2_X4 \u5_seg_h_2/_52_ ( .A1(\u5_seg_h_2/_34_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_10_ ) );
AND2_X1 \u5_seg_h_2/_53_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_10_ ), .ZN(\u5_seg_h_2/_11_ ) );
INV_X1 \u5_seg_h_2/_54_ ( .A(\u5_seg_h_2/_11_ ), .ZN(\u5_seg_h_2/_12_ ) );
INV_X1 \u5_seg_h_2/_55_ ( .A(\u5_seg_h_2/_00_ ), .ZN(\u5_seg_h_2/_13_ ) );
AND2_X4 \u5_seg_h_2/_56_ ( .A1(\u5_seg_h_2/_31_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_14_ ) );
AOI21_X1 \u5_seg_h_2/_57_ ( .A(\u5_seg_h_2/_13_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_15_ ) );
NAND3_X1 \u5_seg_h_2/_58_ ( .A1(\u5_seg_h_2/_07_ ), .A2(\u5_seg_h_2/_12_ ), .A3(\u5_seg_h_2/_15_ ), .ZN(\u5_seg_h_2/_35_ ) );
NAND2_X1 \u5_seg_h_2/_59_ ( .A1(\u5_seg_h_2/_02_ ), .A2(\u5_seg_h_2/_10_ ), .ZN(\u5_seg_h_2/_16_ ) );
AND2_X2 \u5_seg_h_2/_60_ ( .A1(\u5_seg_h_2/_34_ ), .A2(\u5_seg_h_2/_33_ ), .ZN(\u5_seg_h_2/_17_ ) );
NAND2_X1 \u5_seg_h_2/_61_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_17_ ), .ZN(\u5_seg_h_2/_18_ ) );
NAND3_X1 \u5_seg_h_2/_62_ ( .A1(\u5_seg_h_2/_15_ ), .A2(\u5_seg_h_2/_16_ ), .A3(\u5_seg_h_2/_18_ ), .ZN(\u5_seg_h_2/_36_ ) );
NOR3_X1 \u5_seg_h_2/_63_ ( .A1(\u5_seg_h_2/_03_ ), .A2(\u5_seg_h_2/_34_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_19_ ) );
AOI21_X1 \u5_seg_h_2/_64_ ( .A(\u5_seg_h_2/_19_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_20_ ) );
NAND3_X1 \u5_seg_h_2/_65_ ( .A1(\u5_seg_h_2/_05_ ), .A2(\u5_seg_h_2/_03_ ), .A3(\u5_seg_h_2/_31_ ), .ZN(\u5_seg_h_2/_21_ ) );
NAND2_X1 \u5_seg_h_2/_66_ ( .A1(\u5_seg_h_2/_09_ ), .A2(\u5_seg_h_2/_06_ ), .ZN(\u5_seg_h_2/_22_ ) );
NAND4_X1 \u5_seg_h_2/_67_ ( .A1(\u5_seg_h_2/_20_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_21_ ), .A4(\u5_seg_h_2/_22_ ), .ZN(\u5_seg_h_2/_37_ ) );
NAND3_X1 \u5_seg_h_2/_68_ ( .A1(\u5_seg_h_2/_06_ ), .A2(\u5_seg_h_2/_08_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_23_ ) );
AOI22_X1 \u5_seg_h_2/_69_ ( .A1(\u5_seg_h_2/_04_ ), .A2(\u5_seg_h_2/_01_ ), .B1(\u5_seg_h_2/_14_ ), .B2(\u5_seg_h_2/_17_ ), .ZN(\u5_seg_h_2/_24_ ) );
NAND4_X1 \u5_seg_h_2/_70_ ( .A1(\u5_seg_h_2/_12_ ), .A2(\u5_seg_h_2/_15_ ), .A3(\u5_seg_h_2/_23_ ), .A4(\u5_seg_h_2/_24_ ), .ZN(\u5_seg_h_2/_38_ ) );
OAI21_X1 \u5_seg_h_2/_71_ ( .A(\u5_seg_h_2/_17_ ), .B1(\u5_seg_h_2/_08_ ), .B2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_25_ ) );
NAND3_X1 \u5_seg_h_2/_72_ ( .A1(\u5_seg_h_2/_10_ ), .A2(\u5_seg_h_2/_08_ ), .A3(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_26_ ) );
NAND3_X1 \u5_seg_h_2/_73_ ( .A1(\u5_seg_h_2/_25_ ), .A2(\u5_seg_h_2/_26_ ), .A3(\u5_seg_h_2/_00_ ), .ZN(\u5_seg_h_2/_39_ ) );
AND2_X1 \u5_seg_h_2/_74_ ( .A1(\u5_seg_h_2/_08_ ), .A2(\u5_seg_h_2/_32_ ), .ZN(\u5_seg_h_2/_27_ ) );
OAI21_X1 \u5_seg_h_2/_75_ ( .A(\u5_seg_h_2/_04_ ), .B1(\u5_seg_h_2/_27_ ), .B2(\u5_seg_h_2/_09_ ), .ZN(\u5_seg_h_2/_28_ ) );
NAND2_X1 \u5_seg_h_2/_76_ ( .A1(\u5_seg_h_2/_06_ ), .A2(\u5_seg_h_2/_14_ ), .ZN(\u5_seg_h_2/_29_ ) );
NAND4_X1 \u5_seg_h_2/_77_ ( .A1(\u5_seg_h_2/_28_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_25_ ), .A4(\u5_seg_h_2/_29_ ), .ZN(\u5_seg_h_2/_40_ ) );
AOI22_X1 \u5_seg_h_2/_78_ ( .A1(\u5_seg_h_2/_10_ ), .A2(\u5_seg_h_2/_09_ ), .B1(\u5_seg_h_2/_04_ ), .B2(\u5_seg_h_2/_01_ ), .ZN(\u5_seg_h_2/_30_ ) );
NAND4_X1 \u5_seg_h_2/_79_ ( .A1(\u5_seg_h_2/_30_ ), .A2(\u5_seg_h_2/_00_ ), .A3(\u5_seg_h_2/_18_ ), .A4(\u5_seg_h_2/_29_ ), .ZN(\u5_seg_h_2/_41_ ) );
LOGIC1_X1 \u5_seg_h_2/_80_ ( .Z(\u5_seg_h_2/_42_ ) );
BUF_X1 \u5_seg_h_2/_81_ ( .A(\u5_seg_h_2/_42_ ), .Z(\seg_out_0[0] ) );
BUF_X1 \u5_seg_h_2/_82_ ( .A(\key_scan_display[3] ), .Z(\u5_seg_h_2/_34_ ) );
BUF_X1 \u5_seg_h_2/_83_ ( .A(\key_scan_display[2] ), .Z(\u5_seg_h_2/_33_ ) );
BUF_X1 \u5_seg_h_2/_84_ ( .A(\key_scan_display[0] ), .Z(\u5_seg_h_2/_31_ ) );
BUF_X1 \u5_seg_h_2/_85_ ( .A(\key_scan_display[1] ), .Z(\u5_seg_h_2/_32_ ) );
BUF_X1 \u5_seg_h_2/_86_ ( .A(en ), .Z(\u5_seg_h_2/_00_ ) );
BUF_X1 \u5_seg_h_2/_87_ ( .A(\u5_seg_h_2/_35_ ), .Z(\seg_out_0[1] ) );
BUF_X1 \u5_seg_h_2/_88_ ( .A(\u5_seg_h_2/_36_ ), .Z(\seg_out_0[2] ) );
BUF_X1 \u5_seg_h_2/_89_ ( .A(\u5_seg_h_2/_37_ ), .Z(\seg_out_0[3] ) );
BUF_X1 \u5_seg_h_2/_90_ ( .A(\u5_seg_h_2/_38_ ), .Z(\seg_out_0[4] ) );
BUF_X1 \u5_seg_h_2/_91_ ( .A(\u5_seg_h_2/_39_ ), .Z(\seg_out_0[5] ) );
BUF_X1 \u5_seg_h_2/_92_ ( .A(\u5_seg_h_2/_40_ ), .Z(\seg_out_0[6] ) );
BUF_X1 \u5_seg_h_2/_93_ ( .A(\u5_seg_h_2/_41_ ), .Z(\seg_out_0[7] ) );
NOR2_X4 \u6_seg_h_3/_43_ ( .A1(\u6_seg_h_3/_31_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_01_ ) );
INV_X2 \u6_seg_h_3/_44_ ( .A(\u6_seg_h_3/_01_ ), .ZN(\u6_seg_h_3/_02_ ) );
INV_X4 \u6_seg_h_3/_45_ ( .A(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_03_ ) );
NOR2_X2 \u6_seg_h_3/_46_ ( .A1(\u6_seg_h_3/_03_ ), .A2(\u6_seg_h_3/_34_ ), .ZN(\u6_seg_h_3/_04_ ) );
INV_X16 \u6_seg_h_3/_47_ ( .A(\u6_seg_h_3/_34_ ), .ZN(\u6_seg_h_3/_05_ ) );
NOR2_X2 \u6_seg_h_3/_48_ ( .A1(\u6_seg_h_3/_05_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_06_ ) );
OR3_X4 \u6_seg_h_3/_49_ ( .A1(\u6_seg_h_3/_02_ ), .A2(\u6_seg_h_3/_04_ ), .A3(\u6_seg_h_3/_06_ ), .ZN(\u6_seg_h_3/_07_ ) );
INV_X32 \u6_seg_h_3/_50_ ( .A(\u6_seg_h_3/_31_ ), .ZN(\u6_seg_h_3/_08_ ) );
NOR2_X2 \u6_seg_h_3/_51_ ( .A1(\u6_seg_h_3/_08_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_09_ ) );
NOR2_X4 \u6_seg_h_3/_52_ ( .A1(\u6_seg_h_3/_34_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_10_ ) );
AND2_X1 \u6_seg_h_3/_53_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_10_ ), .ZN(\u6_seg_h_3/_11_ ) );
INV_X1 \u6_seg_h_3/_54_ ( .A(\u6_seg_h_3/_11_ ), .ZN(\u6_seg_h_3/_12_ ) );
INV_X1 \u6_seg_h_3/_55_ ( .A(\u6_seg_h_3/_00_ ), .ZN(\u6_seg_h_3/_13_ ) );
AND2_X4 \u6_seg_h_3/_56_ ( .A1(\u6_seg_h_3/_31_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_14_ ) );
AOI21_X1 \u6_seg_h_3/_57_ ( .A(\u6_seg_h_3/_13_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_15_ ) );
NAND3_X1 \u6_seg_h_3/_58_ ( .A1(\u6_seg_h_3/_07_ ), .A2(\u6_seg_h_3/_12_ ), .A3(\u6_seg_h_3/_15_ ), .ZN(\u6_seg_h_3/_35_ ) );
NAND2_X1 \u6_seg_h_3/_59_ ( .A1(\u6_seg_h_3/_02_ ), .A2(\u6_seg_h_3/_10_ ), .ZN(\u6_seg_h_3/_16_ ) );
AND2_X2 \u6_seg_h_3/_60_ ( .A1(\u6_seg_h_3/_34_ ), .A2(\u6_seg_h_3/_33_ ), .ZN(\u6_seg_h_3/_17_ ) );
NAND2_X1 \u6_seg_h_3/_61_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_17_ ), .ZN(\u6_seg_h_3/_18_ ) );
NAND3_X1 \u6_seg_h_3/_62_ ( .A1(\u6_seg_h_3/_15_ ), .A2(\u6_seg_h_3/_16_ ), .A3(\u6_seg_h_3/_18_ ), .ZN(\u6_seg_h_3/_36_ ) );
NOR3_X1 \u6_seg_h_3/_63_ ( .A1(\u6_seg_h_3/_03_ ), .A2(\u6_seg_h_3/_34_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_19_ ) );
AOI21_X1 \u6_seg_h_3/_64_ ( .A(\u6_seg_h_3/_19_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_20_ ) );
NAND3_X1 \u6_seg_h_3/_65_ ( .A1(\u6_seg_h_3/_05_ ), .A2(\u6_seg_h_3/_03_ ), .A3(\u6_seg_h_3/_31_ ), .ZN(\u6_seg_h_3/_21_ ) );
NAND2_X1 \u6_seg_h_3/_66_ ( .A1(\u6_seg_h_3/_09_ ), .A2(\u6_seg_h_3/_06_ ), .ZN(\u6_seg_h_3/_22_ ) );
NAND4_X1 \u6_seg_h_3/_67_ ( .A1(\u6_seg_h_3/_20_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_21_ ), .A4(\u6_seg_h_3/_22_ ), .ZN(\u6_seg_h_3/_37_ ) );
NAND3_X1 \u6_seg_h_3/_68_ ( .A1(\u6_seg_h_3/_06_ ), .A2(\u6_seg_h_3/_08_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_23_ ) );
AOI22_X1 \u6_seg_h_3/_69_ ( .A1(\u6_seg_h_3/_04_ ), .A2(\u6_seg_h_3/_01_ ), .B1(\u6_seg_h_3/_14_ ), .B2(\u6_seg_h_3/_17_ ), .ZN(\u6_seg_h_3/_24_ ) );
NAND4_X1 \u6_seg_h_3/_70_ ( .A1(\u6_seg_h_3/_12_ ), .A2(\u6_seg_h_3/_15_ ), .A3(\u6_seg_h_3/_23_ ), .A4(\u6_seg_h_3/_24_ ), .ZN(\u6_seg_h_3/_38_ ) );
OAI21_X1 \u6_seg_h_3/_71_ ( .A(\u6_seg_h_3/_17_ ), .B1(\u6_seg_h_3/_08_ ), .B2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_25_ ) );
NAND3_X1 \u6_seg_h_3/_72_ ( .A1(\u6_seg_h_3/_10_ ), .A2(\u6_seg_h_3/_08_ ), .A3(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_26_ ) );
NAND3_X1 \u6_seg_h_3/_73_ ( .A1(\u6_seg_h_3/_25_ ), .A2(\u6_seg_h_3/_26_ ), .A3(\u6_seg_h_3/_00_ ), .ZN(\u6_seg_h_3/_39_ ) );
AND2_X1 \u6_seg_h_3/_74_ ( .A1(\u6_seg_h_3/_08_ ), .A2(\u6_seg_h_3/_32_ ), .ZN(\u6_seg_h_3/_27_ ) );
OAI21_X1 \u6_seg_h_3/_75_ ( .A(\u6_seg_h_3/_04_ ), .B1(\u6_seg_h_3/_27_ ), .B2(\u6_seg_h_3/_09_ ), .ZN(\u6_seg_h_3/_28_ ) );
NAND2_X1 \u6_seg_h_3/_76_ ( .A1(\u6_seg_h_3/_06_ ), .A2(\u6_seg_h_3/_14_ ), .ZN(\u6_seg_h_3/_29_ ) );
NAND4_X1 \u6_seg_h_3/_77_ ( .A1(\u6_seg_h_3/_28_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_25_ ), .A4(\u6_seg_h_3/_29_ ), .ZN(\u6_seg_h_3/_40_ ) );
AOI22_X1 \u6_seg_h_3/_78_ ( .A1(\u6_seg_h_3/_10_ ), .A2(\u6_seg_h_3/_09_ ), .B1(\u6_seg_h_3/_04_ ), .B2(\u6_seg_h_3/_01_ ), .ZN(\u6_seg_h_3/_30_ ) );
NAND4_X1 \u6_seg_h_3/_79_ ( .A1(\u6_seg_h_3/_30_ ), .A2(\u6_seg_h_3/_00_ ), .A3(\u6_seg_h_3/_18_ ), .A4(\u6_seg_h_3/_29_ ), .ZN(\u6_seg_h_3/_41_ ) );
LOGIC1_X1 \u6_seg_h_3/_80_ ( .Z(\u6_seg_h_3/_42_ ) );
BUF_X1 \u6_seg_h_3/_81_ ( .A(\u6_seg_h_3/_42_ ), .Z(\seg_out_1[0] ) );
BUF_X1 \u6_seg_h_3/_82_ ( .A(\key_scan_display[7] ), .Z(\u6_seg_h_3/_34_ ) );
BUF_X1 \u6_seg_h_3/_83_ ( .A(\key_scan_display[6] ), .Z(\u6_seg_h_3/_33_ ) );
BUF_X1 \u6_seg_h_3/_84_ ( .A(\key_scan_display[4] ), .Z(\u6_seg_h_3/_31_ ) );
BUF_X1 \u6_seg_h_3/_85_ ( .A(\key_scan_display[5] ), .Z(\u6_seg_h_3/_32_ ) );
BUF_X1 \u6_seg_h_3/_86_ ( .A(en ), .Z(\u6_seg_h_3/_00_ ) );
BUF_X1 \u6_seg_h_3/_87_ ( .A(\u6_seg_h_3/_35_ ), .Z(\seg_out_1[1] ) );
BUF_X1 \u6_seg_h_3/_88_ ( .A(\u6_seg_h_3/_36_ ), .Z(\seg_out_1[2] ) );
BUF_X1 \u6_seg_h_3/_89_ ( .A(\u6_seg_h_3/_37_ ), .Z(\seg_out_1[3] ) );
BUF_X1 \u6_seg_h_3/_90_ ( .A(\u6_seg_h_3/_38_ ), .Z(\seg_out_1[4] ) );
BUF_X1 \u6_seg_h_3/_91_ ( .A(\u6_seg_h_3/_39_ ), .Z(\seg_out_1[5] ) );
BUF_X1 \u6_seg_h_3/_92_ ( .A(\u6_seg_h_3/_40_ ), .Z(\seg_out_1[6] ) );
BUF_X1 \u6_seg_h_3/_93_ ( .A(\u6_seg_h_3/_41_ ), .Z(\seg_out_1[7] ) );
NOR2_X4 \u7_seg_h_4/_43_ ( .A1(\u7_seg_h_4/_31_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_01_ ) );
INV_X2 \u7_seg_h_4/_44_ ( .A(\u7_seg_h_4/_01_ ), .ZN(\u7_seg_h_4/_02_ ) );
INV_X4 \u7_seg_h_4/_45_ ( .A(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_03_ ) );
NOR2_X2 \u7_seg_h_4/_46_ ( .A1(\u7_seg_h_4/_03_ ), .A2(\u7_seg_h_4/_34_ ), .ZN(\u7_seg_h_4/_04_ ) );
INV_X16 \u7_seg_h_4/_47_ ( .A(\u7_seg_h_4/_34_ ), .ZN(\u7_seg_h_4/_05_ ) );
NOR2_X2 \u7_seg_h_4/_48_ ( .A1(\u7_seg_h_4/_05_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_06_ ) );
OR3_X4 \u7_seg_h_4/_49_ ( .A1(\u7_seg_h_4/_02_ ), .A2(\u7_seg_h_4/_04_ ), .A3(\u7_seg_h_4/_06_ ), .ZN(\u7_seg_h_4/_07_ ) );
INV_X32 \u7_seg_h_4/_50_ ( .A(\u7_seg_h_4/_31_ ), .ZN(\u7_seg_h_4/_08_ ) );
NOR2_X2 \u7_seg_h_4/_51_ ( .A1(\u7_seg_h_4/_08_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_09_ ) );
NOR2_X4 \u7_seg_h_4/_52_ ( .A1(\u7_seg_h_4/_34_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_10_ ) );
AND2_X1 \u7_seg_h_4/_53_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_10_ ), .ZN(\u7_seg_h_4/_11_ ) );
INV_X1 \u7_seg_h_4/_54_ ( .A(\u7_seg_h_4/_11_ ), .ZN(\u7_seg_h_4/_12_ ) );
INV_X1 \u7_seg_h_4/_55_ ( .A(\u7_seg_h_4/_00_ ), .ZN(\u7_seg_h_4/_13_ ) );
AND2_X4 \u7_seg_h_4/_56_ ( .A1(\u7_seg_h_4/_31_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_14_ ) );
AOI21_X1 \u7_seg_h_4/_57_ ( .A(\u7_seg_h_4/_13_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_15_ ) );
NAND3_X1 \u7_seg_h_4/_58_ ( .A1(\u7_seg_h_4/_07_ ), .A2(\u7_seg_h_4/_12_ ), .A3(\u7_seg_h_4/_15_ ), .ZN(\u7_seg_h_4/_35_ ) );
NAND2_X1 \u7_seg_h_4/_59_ ( .A1(\u7_seg_h_4/_02_ ), .A2(\u7_seg_h_4/_10_ ), .ZN(\u7_seg_h_4/_16_ ) );
AND2_X2 \u7_seg_h_4/_60_ ( .A1(\u7_seg_h_4/_34_ ), .A2(\u7_seg_h_4/_33_ ), .ZN(\u7_seg_h_4/_17_ ) );
NAND2_X1 \u7_seg_h_4/_61_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_17_ ), .ZN(\u7_seg_h_4/_18_ ) );
NAND3_X1 \u7_seg_h_4/_62_ ( .A1(\u7_seg_h_4/_15_ ), .A2(\u7_seg_h_4/_16_ ), .A3(\u7_seg_h_4/_18_ ), .ZN(\u7_seg_h_4/_36_ ) );
NOR3_X1 \u7_seg_h_4/_63_ ( .A1(\u7_seg_h_4/_03_ ), .A2(\u7_seg_h_4/_34_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_19_ ) );
AOI21_X1 \u7_seg_h_4/_64_ ( .A(\u7_seg_h_4/_19_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_20_ ) );
NAND3_X1 \u7_seg_h_4/_65_ ( .A1(\u7_seg_h_4/_05_ ), .A2(\u7_seg_h_4/_03_ ), .A3(\u7_seg_h_4/_31_ ), .ZN(\u7_seg_h_4/_21_ ) );
NAND2_X1 \u7_seg_h_4/_66_ ( .A1(\u7_seg_h_4/_09_ ), .A2(\u7_seg_h_4/_06_ ), .ZN(\u7_seg_h_4/_22_ ) );
NAND4_X1 \u7_seg_h_4/_67_ ( .A1(\u7_seg_h_4/_20_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_21_ ), .A4(\u7_seg_h_4/_22_ ), .ZN(\u7_seg_h_4/_37_ ) );
NAND3_X1 \u7_seg_h_4/_68_ ( .A1(\u7_seg_h_4/_06_ ), .A2(\u7_seg_h_4/_08_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_23_ ) );
AOI22_X1 \u7_seg_h_4/_69_ ( .A1(\u7_seg_h_4/_04_ ), .A2(\u7_seg_h_4/_01_ ), .B1(\u7_seg_h_4/_14_ ), .B2(\u7_seg_h_4/_17_ ), .ZN(\u7_seg_h_4/_24_ ) );
NAND4_X1 \u7_seg_h_4/_70_ ( .A1(\u7_seg_h_4/_12_ ), .A2(\u7_seg_h_4/_15_ ), .A3(\u7_seg_h_4/_23_ ), .A4(\u7_seg_h_4/_24_ ), .ZN(\u7_seg_h_4/_38_ ) );
OAI21_X1 \u7_seg_h_4/_71_ ( .A(\u7_seg_h_4/_17_ ), .B1(\u7_seg_h_4/_08_ ), .B2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_25_ ) );
NAND3_X1 \u7_seg_h_4/_72_ ( .A1(\u7_seg_h_4/_10_ ), .A2(\u7_seg_h_4/_08_ ), .A3(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_26_ ) );
NAND3_X1 \u7_seg_h_4/_73_ ( .A1(\u7_seg_h_4/_25_ ), .A2(\u7_seg_h_4/_26_ ), .A3(\u7_seg_h_4/_00_ ), .ZN(\u7_seg_h_4/_39_ ) );
AND2_X1 \u7_seg_h_4/_74_ ( .A1(\u7_seg_h_4/_08_ ), .A2(\u7_seg_h_4/_32_ ), .ZN(\u7_seg_h_4/_27_ ) );
OAI21_X1 \u7_seg_h_4/_75_ ( .A(\u7_seg_h_4/_04_ ), .B1(\u7_seg_h_4/_27_ ), .B2(\u7_seg_h_4/_09_ ), .ZN(\u7_seg_h_4/_28_ ) );
NAND2_X1 \u7_seg_h_4/_76_ ( .A1(\u7_seg_h_4/_06_ ), .A2(\u7_seg_h_4/_14_ ), .ZN(\u7_seg_h_4/_29_ ) );
NAND4_X1 \u7_seg_h_4/_77_ ( .A1(\u7_seg_h_4/_28_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_25_ ), .A4(\u7_seg_h_4/_29_ ), .ZN(\u7_seg_h_4/_40_ ) );
AOI22_X1 \u7_seg_h_4/_78_ ( .A1(\u7_seg_h_4/_10_ ), .A2(\u7_seg_h_4/_09_ ), .B1(\u7_seg_h_4/_04_ ), .B2(\u7_seg_h_4/_01_ ), .ZN(\u7_seg_h_4/_30_ ) );
NAND4_X1 \u7_seg_h_4/_79_ ( .A1(\u7_seg_h_4/_30_ ), .A2(\u7_seg_h_4/_00_ ), .A3(\u7_seg_h_4/_18_ ), .A4(\u7_seg_h_4/_29_ ), .ZN(\u7_seg_h_4/_41_ ) );
LOGIC1_X1 \u7_seg_h_4/_80_ ( .Z(\u7_seg_h_4/_42_ ) );
BUF_X1 \u7_seg_h_4/_81_ ( .A(\u7_seg_h_4/_42_ ), .Z(\seg_out_4[0] ) );
BUF_X1 \u7_seg_h_4/_82_ ( .A(\high_units[3] ), .Z(\u7_seg_h_4/_34_ ) );
BUF_X1 \u7_seg_h_4/_83_ ( .A(\high_units[2] ), .Z(\u7_seg_h_4/_33_ ) );
BUF_X1 \u7_seg_h_4/_84_ ( .A(\high_units[0] ), .Z(\u7_seg_h_4/_31_ ) );
BUF_X1 \u7_seg_h_4/_85_ ( .A(\high_units[1] ), .Z(\u7_seg_h_4/_32_ ) );
BUF_X1 \u7_seg_h_4/_86_ ( .A(_132_ ), .Z(\u7_seg_h_4/_00_ ) );
BUF_X1 \u7_seg_h_4/_87_ ( .A(\u7_seg_h_4/_35_ ), .Z(\seg_out_4[1] ) );
BUF_X1 \u7_seg_h_4/_88_ ( .A(\u7_seg_h_4/_36_ ), .Z(\seg_out_4[2] ) );
BUF_X1 \u7_seg_h_4/_89_ ( .A(\u7_seg_h_4/_37_ ), .Z(\seg_out_4[3] ) );
BUF_X1 \u7_seg_h_4/_90_ ( .A(\u7_seg_h_4/_38_ ), .Z(\seg_out_4[4] ) );
BUF_X1 \u7_seg_h_4/_91_ ( .A(\u7_seg_h_4/_39_ ), .Z(\seg_out_4[5] ) );
BUF_X1 \u7_seg_h_4/_92_ ( .A(\u7_seg_h_4/_40_ ), .Z(\seg_out_4[6] ) );
BUF_X1 \u7_seg_h_4/_93_ ( .A(\u7_seg_h_4/_41_ ), .Z(\seg_out_4[7] ) );
NOR2_X4 \u8_seg_h_5/_43_ ( .A1(\u8_seg_h_5/_31_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_01_ ) );
INV_X2 \u8_seg_h_5/_44_ ( .A(\u8_seg_h_5/_01_ ), .ZN(\u8_seg_h_5/_02_ ) );
INV_X4 \u8_seg_h_5/_45_ ( .A(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_03_ ) );
NOR2_X2 \u8_seg_h_5/_46_ ( .A1(\u8_seg_h_5/_03_ ), .A2(\u8_seg_h_5/_34_ ), .ZN(\u8_seg_h_5/_04_ ) );
INV_X16 \u8_seg_h_5/_47_ ( .A(\u8_seg_h_5/_34_ ), .ZN(\u8_seg_h_5/_05_ ) );
NOR2_X2 \u8_seg_h_5/_48_ ( .A1(\u8_seg_h_5/_05_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_06_ ) );
OR3_X4 \u8_seg_h_5/_49_ ( .A1(\u8_seg_h_5/_02_ ), .A2(\u8_seg_h_5/_04_ ), .A3(\u8_seg_h_5/_06_ ), .ZN(\u8_seg_h_5/_07_ ) );
INV_X32 \u8_seg_h_5/_50_ ( .A(\u8_seg_h_5/_31_ ), .ZN(\u8_seg_h_5/_08_ ) );
NOR2_X2 \u8_seg_h_5/_51_ ( .A1(\u8_seg_h_5/_08_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_09_ ) );
NOR2_X4 \u8_seg_h_5/_52_ ( .A1(\u8_seg_h_5/_34_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_10_ ) );
AND2_X1 \u8_seg_h_5/_53_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_10_ ), .ZN(\u8_seg_h_5/_11_ ) );
INV_X1 \u8_seg_h_5/_54_ ( .A(\u8_seg_h_5/_11_ ), .ZN(\u8_seg_h_5/_12_ ) );
INV_X1 \u8_seg_h_5/_55_ ( .A(\u8_seg_h_5/_00_ ), .ZN(\u8_seg_h_5/_13_ ) );
AND2_X4 \u8_seg_h_5/_56_ ( .A1(\u8_seg_h_5/_31_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_14_ ) );
AOI21_X1 \u8_seg_h_5/_57_ ( .A(\u8_seg_h_5/_13_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_15_ ) );
NAND3_X1 \u8_seg_h_5/_58_ ( .A1(\u8_seg_h_5/_07_ ), .A2(\u8_seg_h_5/_12_ ), .A3(\u8_seg_h_5/_15_ ), .ZN(\u8_seg_h_5/_35_ ) );
NAND2_X1 \u8_seg_h_5/_59_ ( .A1(\u8_seg_h_5/_02_ ), .A2(\u8_seg_h_5/_10_ ), .ZN(\u8_seg_h_5/_16_ ) );
AND2_X2 \u8_seg_h_5/_60_ ( .A1(\u8_seg_h_5/_34_ ), .A2(\u8_seg_h_5/_33_ ), .ZN(\u8_seg_h_5/_17_ ) );
NAND2_X1 \u8_seg_h_5/_61_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_17_ ), .ZN(\u8_seg_h_5/_18_ ) );
NAND3_X1 \u8_seg_h_5/_62_ ( .A1(\u8_seg_h_5/_15_ ), .A2(\u8_seg_h_5/_16_ ), .A3(\u8_seg_h_5/_18_ ), .ZN(\u8_seg_h_5/_36_ ) );
NOR3_X1 \u8_seg_h_5/_63_ ( .A1(\u8_seg_h_5/_03_ ), .A2(\u8_seg_h_5/_34_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_19_ ) );
AOI21_X1 \u8_seg_h_5/_64_ ( .A(\u8_seg_h_5/_19_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_20_ ) );
NAND3_X1 \u8_seg_h_5/_65_ ( .A1(\u8_seg_h_5/_05_ ), .A2(\u8_seg_h_5/_03_ ), .A3(\u8_seg_h_5/_31_ ), .ZN(\u8_seg_h_5/_21_ ) );
NAND2_X1 \u8_seg_h_5/_66_ ( .A1(\u8_seg_h_5/_09_ ), .A2(\u8_seg_h_5/_06_ ), .ZN(\u8_seg_h_5/_22_ ) );
NAND4_X1 \u8_seg_h_5/_67_ ( .A1(\u8_seg_h_5/_20_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_21_ ), .A4(\u8_seg_h_5/_22_ ), .ZN(\u8_seg_h_5/_37_ ) );
NAND3_X1 \u8_seg_h_5/_68_ ( .A1(\u8_seg_h_5/_06_ ), .A2(\u8_seg_h_5/_08_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_23_ ) );
AOI22_X1 \u8_seg_h_5/_69_ ( .A1(\u8_seg_h_5/_04_ ), .A2(\u8_seg_h_5/_01_ ), .B1(\u8_seg_h_5/_14_ ), .B2(\u8_seg_h_5/_17_ ), .ZN(\u8_seg_h_5/_24_ ) );
NAND4_X1 \u8_seg_h_5/_70_ ( .A1(\u8_seg_h_5/_12_ ), .A2(\u8_seg_h_5/_15_ ), .A3(\u8_seg_h_5/_23_ ), .A4(\u8_seg_h_5/_24_ ), .ZN(\u8_seg_h_5/_38_ ) );
OAI21_X1 \u8_seg_h_5/_71_ ( .A(\u8_seg_h_5/_17_ ), .B1(\u8_seg_h_5/_08_ ), .B2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_25_ ) );
NAND3_X1 \u8_seg_h_5/_72_ ( .A1(\u8_seg_h_5/_10_ ), .A2(\u8_seg_h_5/_08_ ), .A3(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_26_ ) );
NAND3_X1 \u8_seg_h_5/_73_ ( .A1(\u8_seg_h_5/_25_ ), .A2(\u8_seg_h_5/_26_ ), .A3(\u8_seg_h_5/_00_ ), .ZN(\u8_seg_h_5/_39_ ) );
AND2_X1 \u8_seg_h_5/_74_ ( .A1(\u8_seg_h_5/_08_ ), .A2(\u8_seg_h_5/_32_ ), .ZN(\u8_seg_h_5/_27_ ) );
OAI21_X1 \u8_seg_h_5/_75_ ( .A(\u8_seg_h_5/_04_ ), .B1(\u8_seg_h_5/_27_ ), .B2(\u8_seg_h_5/_09_ ), .ZN(\u8_seg_h_5/_28_ ) );
NAND2_X1 \u8_seg_h_5/_76_ ( .A1(\u8_seg_h_5/_06_ ), .A2(\u8_seg_h_5/_14_ ), .ZN(\u8_seg_h_5/_29_ ) );
NAND4_X1 \u8_seg_h_5/_77_ ( .A1(\u8_seg_h_5/_28_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_25_ ), .A4(\u8_seg_h_5/_29_ ), .ZN(\u8_seg_h_5/_40_ ) );
AOI22_X1 \u8_seg_h_5/_78_ ( .A1(\u8_seg_h_5/_10_ ), .A2(\u8_seg_h_5/_09_ ), .B1(\u8_seg_h_5/_04_ ), .B2(\u8_seg_h_5/_01_ ), .ZN(\u8_seg_h_5/_30_ ) );
NAND4_X1 \u8_seg_h_5/_79_ ( .A1(\u8_seg_h_5/_30_ ), .A2(\u8_seg_h_5/_00_ ), .A3(\u8_seg_h_5/_18_ ), .A4(\u8_seg_h_5/_29_ ), .ZN(\u8_seg_h_5/_41_ ) );
LOGIC1_X1 \u8_seg_h_5/_80_ ( .Z(\u8_seg_h_5/_42_ ) );
BUF_X1 \u8_seg_h_5/_81_ ( .A(\u8_seg_h_5/_42_ ), .Z(\seg_out_5[0] ) );
BUF_X1 \u8_seg_h_5/_82_ ( .A(\high_tens[3] ), .Z(\u8_seg_h_5/_34_ ) );
BUF_X1 \u8_seg_h_5/_83_ ( .A(\high_tens[2] ), .Z(\u8_seg_h_5/_33_ ) );
BUF_X1 \u8_seg_h_5/_84_ ( .A(\high_tens[0] ), .Z(\u8_seg_h_5/_31_ ) );
BUF_X1 \u8_seg_h_5/_85_ ( .A(\high_tens[1] ), .Z(\u8_seg_h_5/_32_ ) );
BUF_X1 \u8_seg_h_5/_86_ ( .A(_132_ ), .Z(\u8_seg_h_5/_00_ ) );
BUF_X1 \u8_seg_h_5/_87_ ( .A(\u8_seg_h_5/_35_ ), .Z(\seg_out_5[1] ) );
BUF_X1 \u8_seg_h_5/_88_ ( .A(\u8_seg_h_5/_36_ ), .Z(\seg_out_5[2] ) );
BUF_X1 \u8_seg_h_5/_89_ ( .A(\u8_seg_h_5/_37_ ), .Z(\seg_out_5[3] ) );
BUF_X1 \u8_seg_h_5/_90_ ( .A(\u8_seg_h_5/_38_ ), .Z(\seg_out_5[4] ) );
BUF_X1 \u8_seg_h_5/_91_ ( .A(\u8_seg_h_5/_39_ ), .Z(\seg_out_5[5] ) );
BUF_X1 \u8_seg_h_5/_92_ ( .A(\u8_seg_h_5/_40_ ), .Z(\seg_out_5[6] ) );
BUF_X1 \u8_seg_h_5/_93_ ( .A(\u8_seg_h_5/_41_ ), .Z(\seg_out_5[7] ) );
BUF_X8 fanout_buf_1 ( .A(\u0_ps2_kb/_0476_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(clrn ), .Z(fanout_net_2 ) );

endmodule
